magic
tech sky130A
magscale 1 2
timestamp 1655908342
<< viali >>
rect 41061 57409 41095 57443
rect 41705 57341 41739 57375
rect 7849 56797 7883 56831
rect 9045 56797 9079 56831
rect 26065 56797 26099 56831
rect 33609 56797 33643 56831
rect 35725 56797 35759 56831
rect 42533 56797 42567 56831
rect 43177 56797 43211 56831
rect 50169 56797 50203 56831
rect 52929 56797 52963 56831
rect 43269 56389 43303 56423
rect 8493 56321 8527 56355
rect 8953 56321 8987 56355
rect 33517 56321 33551 56355
rect 49893 56321 49927 56355
rect 52837 56321 52871 56355
rect 7757 56253 7791 56287
rect 8309 56253 8343 56287
rect 9137 56253 9171 56287
rect 9689 56253 9723 56287
rect 33701 56253 33735 56287
rect 34161 56253 34195 56287
rect 44925 56253 44959 56287
rect 45109 56253 45143 56287
rect 50077 56253 50111 56287
rect 51089 56253 51123 56287
rect 53021 56253 53055 56287
rect 53297 56253 53331 56287
rect 42625 56117 42659 56151
rect 33701 55913 33735 55947
rect 44373 55913 44407 55947
rect 50261 55913 50295 55947
rect 53205 55913 53239 55947
rect 25973 55777 26007 55811
rect 26433 55777 26467 55811
rect 35725 55777 35759 55811
rect 36185 55777 36219 55811
rect 41981 55777 42015 55811
rect 42444 55777 42478 55811
rect 33609 55709 33643 55743
rect 42717 55709 42751 55743
rect 44465 55709 44499 55743
rect 50361 55711 50395 55745
rect 53297 55709 53331 55743
rect 26157 55641 26191 55675
rect 35909 55641 35943 55675
rect 42447 55573 42481 55607
rect 43821 55573 43855 55607
rect 9137 55369 9171 55403
rect 26157 55369 26191 55403
rect 35909 55369 35943 55403
rect 42441 55369 42475 55403
rect 43814 55369 43848 55403
rect 9045 55233 9079 55267
rect 26065 55233 26099 55267
rect 35817 55233 35851 55267
rect 43545 55233 43579 55267
rect 44281 55233 44315 55267
rect 43818 55165 43852 55199
rect 44189 54825 44223 54859
rect 42349 54689 42383 54723
rect 42855 54689 42889 54723
rect 2053 54621 2087 54655
rect 43085 54621 43119 54655
rect 42815 54485 42849 54519
rect 1961 54145 1995 54179
rect 46305 54145 46339 54179
rect 46489 54145 46523 54179
rect 2145 54077 2179 54111
rect 2789 54077 2823 54111
rect 46305 53941 46339 53975
rect 2421 53737 2455 53771
rect 46765 53737 46799 53771
rect 45477 53669 45511 53703
rect 2513 53533 2547 53567
rect 42625 53533 42659 53567
rect 45753 53533 45787 53567
rect 46581 53533 46615 53567
rect 45477 53465 45511 53499
rect 45661 53397 45695 53431
rect 44281 53193 44315 53227
rect 46590 53125 46624 53159
rect 49801 53125 49835 53159
rect 42441 53057 42475 53091
rect 42764 53057 42798 53091
rect 48053 53057 48087 53091
rect 49065 53057 49099 53091
rect 42904 52989 42938 53023
rect 43177 52989 43211 53023
rect 46857 52989 46891 53023
rect 47777 52989 47811 53023
rect 50261 52989 50295 53023
rect 50353 52989 50387 53023
rect 47961 52921 47995 52955
rect 49801 52921 49835 52955
rect 45477 52853 45511 52887
rect 47869 52853 47903 52887
rect 49249 52853 49283 52887
rect 50537 52853 50571 52887
rect 41429 52649 41463 52683
rect 43729 52649 43763 52683
rect 46857 52649 46891 52683
rect 49341 52649 49375 52683
rect 46397 52581 46431 52615
rect 48881 52581 48915 52615
rect 50261 52581 50295 52615
rect 41889 52513 41923 52547
rect 42395 52513 42429 52547
rect 44189 52513 44223 52547
rect 45017 52513 45051 52547
rect 50813 52513 50847 52547
rect 42625 52445 42659 52479
rect 45284 52445 45318 52479
rect 47041 52445 47075 52479
rect 47501 52445 47535 52479
rect 47768 52445 47802 52479
rect 49341 52445 49375 52479
rect 49617 52445 49651 52479
rect 50721 52445 50755 52479
rect 49525 52377 49559 52411
rect 50261 52377 50295 52411
rect 42355 52309 42389 52343
rect 50997 52309 51031 52343
rect 42441 52105 42475 52139
rect 43814 52105 43848 52139
rect 45569 52105 45603 52139
rect 46489 52105 46523 52139
rect 47961 52105 47995 52139
rect 49525 52105 49559 52139
rect 47593 52037 47627 52071
rect 47809 52037 47843 52071
rect 49985 52037 50019 52071
rect 46029 51969 46063 52003
rect 46949 51969 46983 52003
rect 49433 51969 49467 52003
rect 51067 51975 51101 52009
rect 51549 51969 51583 52003
rect 43545 51901 43579 51935
rect 43775 51901 43809 51935
rect 44281 51901 44315 51935
rect 50813 51901 50847 51935
rect 49985 51833 50019 51867
rect 45937 51765 45971 51799
rect 46673 51765 46707 51799
rect 47777 51765 47811 51799
rect 49249 51765 49283 51799
rect 50537 51765 50571 51799
rect 50721 51765 50755 51799
rect 51733 51765 51767 51799
rect 46029 51561 46063 51595
rect 47409 51425 47443 51459
rect 45017 51357 45051 51391
rect 45201 51357 45235 51391
rect 46213 51357 46247 51391
rect 46397 51357 46431 51391
rect 47593 51357 47627 51391
rect 50629 51357 50663 51391
rect 47777 51289 47811 51323
rect 45109 51221 45143 51255
rect 50813 51221 50847 51255
rect 48605 51017 48639 51051
rect 44741 50881 44775 50915
rect 44925 50881 44959 50915
rect 45845 50881 45879 50915
rect 46029 50881 46063 50915
rect 48421 50881 48455 50915
rect 49433 50881 49467 50915
rect 50445 50881 50479 50915
rect 44741 50677 44775 50711
rect 46029 50677 46063 50711
rect 49249 50677 49283 50711
rect 50353 50677 50387 50711
rect 48789 50405 48823 50439
rect 48605 50337 48639 50371
rect 37565 50269 37599 50303
rect 47685 50269 47719 50303
rect 47961 50269 47995 50303
rect 48145 50269 48179 50303
rect 37832 50201 37866 50235
rect 49065 50201 49099 50235
rect 38945 50133 38979 50167
rect 47501 50133 47535 50167
rect 37933 49929 37967 49963
rect 43735 49929 43769 49963
rect 50819 49929 50853 49963
rect 52193 49929 52227 49963
rect 47838 49861 47872 49895
rect 38117 49793 38151 49827
rect 38393 49793 38427 49827
rect 38577 49793 38611 49827
rect 39497 49793 39531 49827
rect 40509 49793 40543 49827
rect 40776 49793 40810 49827
rect 43269 49793 43303 49827
rect 1961 49725 1995 49759
rect 2145 49725 2179 49759
rect 2789 49725 2823 49759
rect 39681 49725 39715 49759
rect 43732 49725 43766 49759
rect 44005 49725 44039 49759
rect 47593 49725 47627 49759
rect 50353 49725 50387 49759
rect 50816 49725 50850 49759
rect 51089 49725 51123 49759
rect 39313 49589 39347 49623
rect 41889 49589 41923 49623
rect 45109 49589 45143 49623
rect 48973 49589 49007 49623
rect 2053 49385 2087 49419
rect 52009 49385 52043 49419
rect 54309 49385 54343 49419
rect 39221 49317 39255 49351
rect 39865 49317 39899 49351
rect 36277 49249 36311 49283
rect 40141 49249 40175 49283
rect 41340 49249 41374 49283
rect 45480 49249 45514 49283
rect 48240 49249 48274 49283
rect 48513 49249 48547 49283
rect 50632 49249 50666 49283
rect 52792 49249 52826 49283
rect 52932 49249 52966 49283
rect 53205 49249 53239 49283
rect 40049 49181 40083 49215
rect 40233 49181 40267 49215
rect 40325 49181 40359 49215
rect 40877 49181 40911 49215
rect 41613 49181 41647 49215
rect 45017 49181 45051 49215
rect 45753 49181 45787 49215
rect 47777 49181 47811 49215
rect 50169 49181 50203 49215
rect 50905 49181 50939 49215
rect 52469 49181 52503 49215
rect 36544 49113 36578 49147
rect 38853 49113 38887 49147
rect 37657 49045 37691 49079
rect 39313 49045 39347 49079
rect 41343 49045 41377 49079
rect 42717 49045 42751 49079
rect 45483 49045 45517 49079
rect 46857 49045 46891 49079
rect 48243 49045 48277 49079
rect 49617 49045 49651 49079
rect 50635 49045 50669 49079
rect 2421 48841 2455 48875
rect 36737 48841 36771 48875
rect 37565 48841 37599 48875
rect 38393 48841 38427 48875
rect 39405 48841 39439 48875
rect 39773 48841 39807 48875
rect 40693 48841 40727 48875
rect 42907 48841 42941 48875
rect 44281 48841 44315 48875
rect 45753 48841 45787 48875
rect 49071 48841 49105 48875
rect 50445 48841 50479 48875
rect 37733 48773 37767 48807
rect 37933 48773 37967 48807
rect 47685 48773 47719 48807
rect 2513 48705 2547 48739
rect 36737 48705 36771 48739
rect 38669 48705 38703 48739
rect 38761 48705 38795 48739
rect 39681 48705 39715 48739
rect 40509 48705 40543 48739
rect 42441 48705 42475 48739
rect 43177 48705 43211 48739
rect 45017 48705 45051 48739
rect 36461 48637 36495 48671
rect 38577 48637 38611 48671
rect 38853 48637 38887 48671
rect 39589 48637 39623 48671
rect 39957 48637 39991 48671
rect 40049 48637 40083 48671
rect 42904 48637 42938 48671
rect 44741 48637 44775 48671
rect 48605 48637 48639 48671
rect 49111 48637 49145 48671
rect 49341 48637 49375 48671
rect 36645 48569 36679 48603
rect 48053 48569 48087 48603
rect 37749 48501 37783 48535
rect 48145 48501 48179 48535
rect 37473 48297 37507 48331
rect 48237 48297 48271 48331
rect 47593 48229 47627 48263
rect 40141 48161 40175 48195
rect 45753 48161 45787 48195
rect 46216 48161 46250 48195
rect 46489 48161 46523 48195
rect 2053 48093 2087 48127
rect 37197 48093 37231 48127
rect 39865 48093 39899 48127
rect 48421 48093 48455 48127
rect 37473 48025 37507 48059
rect 37289 47957 37323 47991
rect 46219 47957 46253 47991
rect 40515 47753 40549 47787
rect 41889 47753 41923 47787
rect 45661 47753 45695 47787
rect 36645 47685 36679 47719
rect 1961 47617 1995 47651
rect 36369 47617 36403 47651
rect 36737 47617 36771 47651
rect 37749 47617 37783 47651
rect 46397 47617 46431 47651
rect 46673 47617 46707 47651
rect 2145 47549 2179 47583
rect 2789 47549 2823 47583
rect 37473 47549 37507 47583
rect 40049 47549 40083 47583
rect 40512 47549 40546 47583
rect 40785 47549 40819 47583
rect 36369 47413 36403 47447
rect 36461 47413 36495 47447
rect 2421 47209 2455 47243
rect 38209 47209 38243 47243
rect 39313 47209 39347 47243
rect 51825 47209 51859 47243
rect 57989 47141 58023 47175
rect 38945 47073 38979 47107
rect 40141 47073 40175 47107
rect 43453 47073 43487 47107
rect 50813 47073 50847 47107
rect 52285 47073 52319 47107
rect 52608 47073 52642 47107
rect 52791 47073 52825 47107
rect 53021 47073 53055 47107
rect 2513 47005 2547 47039
rect 36369 47005 36403 47039
rect 36625 47005 36659 47039
rect 38393 47005 38427 47039
rect 38485 47005 38519 47039
rect 39129 47005 39163 47039
rect 39865 47005 39899 47039
rect 42993 47005 43027 47039
rect 43729 47005 43763 47039
rect 51089 47005 51123 47039
rect 58173 47005 58207 47039
rect 38209 46937 38243 46971
rect 37749 46869 37783 46903
rect 44465 46869 44499 46903
rect 54125 46869 54159 46903
rect 40515 46665 40549 46699
rect 41889 46665 41923 46699
rect 44465 46665 44499 46699
rect 48966 46665 49000 46699
rect 52745 46665 52779 46699
rect 37381 46597 37415 46631
rect 52929 46597 52963 46631
rect 37289 46529 37323 46563
rect 37565 46529 37599 46563
rect 42948 46529 42982 46563
rect 48697 46529 48731 46563
rect 51181 46529 51215 46563
rect 40049 46461 40083 46495
rect 40512 46479 40546 46513
rect 40785 46461 40819 46495
rect 42625 46461 42659 46495
rect 43088 46461 43122 46495
rect 43361 46461 43395 46495
rect 48927 46461 48961 46495
rect 49433 46461 49467 46495
rect 47593 46393 47627 46427
rect 53297 46393 53331 46427
rect 37565 46325 37599 46359
rect 50997 46325 51031 46359
rect 52929 46325 52963 46359
rect 52101 46053 52135 46087
rect 36277 45985 36311 46019
rect 38117 45985 38151 46019
rect 44465 45985 44499 46019
rect 47777 45985 47811 46019
rect 48100 45985 48134 46019
rect 48240 45985 48274 46019
rect 53021 45985 53055 46019
rect 38393 45917 38427 45951
rect 44189 45917 44223 45951
rect 45661 45917 45695 45951
rect 48513 45917 48547 45951
rect 51089 45917 51123 45951
rect 51365 45917 51399 45951
rect 52745 45917 52779 45951
rect 36544 45849 36578 45883
rect 45928 45849 45962 45883
rect 37657 45781 37691 45815
rect 43453 45781 43487 45815
rect 47041 45781 47075 45815
rect 49617 45781 49651 45815
rect 40423 45577 40457 45611
rect 41797 45577 41831 45611
rect 48973 45577 49007 45611
rect 50346 45577 50380 45611
rect 52745 45577 52779 45611
rect 52929 45577 52963 45611
rect 37289 45509 37323 45543
rect 46857 45509 46891 45543
rect 37473 45441 37507 45475
rect 37749 45441 37783 45475
rect 44373 45441 44407 45475
rect 45109 45441 45143 45475
rect 45569 45441 45603 45475
rect 45845 45441 45879 45475
rect 46489 45441 46523 45475
rect 46949 45441 46983 45475
rect 50077 45441 50111 45475
rect 53297 45441 53331 45475
rect 39957 45373 39991 45407
rect 40420 45391 40454 45425
rect 40693 45373 40727 45407
rect 45477 45373 45511 45407
rect 50307 45373 50341 45407
rect 50813 45373 50847 45407
rect 2053 45237 2087 45271
rect 37657 45237 37691 45271
rect 43913 45237 43947 45271
rect 44281 45237 44315 45271
rect 46627 45237 46661 45271
rect 46765 45237 46799 45271
rect 52929 45237 52963 45271
rect 41705 45033 41739 45067
rect 45845 45033 45879 45067
rect 46949 45033 46983 45067
rect 47409 45033 47443 45067
rect 47593 45033 47627 45067
rect 36921 44965 36955 44999
rect 37749 44965 37783 44999
rect 36737 44897 36771 44931
rect 40328 44897 40362 44931
rect 50445 44897 50479 44931
rect 51917 44897 51951 44931
rect 2513 44829 2547 44863
rect 37013 44829 37047 44863
rect 37473 44829 37507 44863
rect 37749 44829 37783 44863
rect 39865 44829 39899 44863
rect 40601 44829 40635 44863
rect 43085 44829 43119 44863
rect 45385 44829 45419 44863
rect 45661 44829 45695 44863
rect 46305 44829 46339 44863
rect 46489 44829 46523 44863
rect 46581 44829 46615 44863
rect 46719 44829 46753 44863
rect 47593 44829 47627 44863
rect 47685 44829 47719 44863
rect 48053 44829 48087 44863
rect 50721 44829 50755 44863
rect 52193 44829 52227 44863
rect 43352 44761 43386 44795
rect 45477 44761 45511 44795
rect 2421 44693 2455 44727
rect 37013 44693 37047 44727
rect 37565 44693 37599 44727
rect 40331 44693 40365 44727
rect 44465 44693 44499 44727
rect 51457 44693 51491 44727
rect 52929 44693 52963 44727
rect 38669 44489 38703 44523
rect 39513 44489 39547 44523
rect 39681 44489 39715 44523
rect 40141 44489 40175 44523
rect 43729 44489 43763 44523
rect 49623 44489 49657 44523
rect 53021 44489 53055 44523
rect 2145 44421 2179 44455
rect 37534 44421 37568 44455
rect 39313 44421 39347 44455
rect 52745 44421 52779 44455
rect 1961 44353 1995 44387
rect 37289 44353 37323 44387
rect 40877 44353 40911 44387
rect 43913 44353 43947 44387
rect 44649 44353 44683 44387
rect 46213 44353 46247 44387
rect 46305 44353 46339 44387
rect 46489 44353 46523 44387
rect 49893 44353 49927 44387
rect 53021 44353 53055 44387
rect 2789 44285 2823 44319
rect 41153 44285 41187 44319
rect 44925 44285 44959 44319
rect 49157 44285 49191 44319
rect 49663 44285 49697 44319
rect 52929 44285 52963 44319
rect 46489 44217 46523 44251
rect 39497 44149 39531 44183
rect 50997 44149 51031 44183
rect 40509 43945 40543 43979
rect 46673 43945 46707 43979
rect 38025 43877 38059 43911
rect 41521 43809 41555 43843
rect 37289 43741 37323 43775
rect 37473 43741 37507 43775
rect 37565 43741 37599 43775
rect 38301 43741 38335 43775
rect 41245 43741 41279 43775
rect 44097 43741 44131 43775
rect 44281 43741 44315 43775
rect 46765 43741 46799 43775
rect 38025 43673 38059 43707
rect 37105 43605 37139 43639
rect 38209 43605 38243 43639
rect 44281 43605 44315 43639
rect 40331 43401 40365 43435
rect 41705 43401 41739 43435
rect 46121 43401 46155 43435
rect 49610 43401 49644 43435
rect 53205 43401 53239 43435
rect 36645 43333 36679 43367
rect 37534 43333 37568 43367
rect 43913 43333 43947 43367
rect 46581 43333 46615 43367
rect 36553 43265 36587 43299
rect 36737 43265 36771 43299
rect 44097 43265 44131 43299
rect 45293 43265 45327 43299
rect 46305 43265 46339 43299
rect 52745 43265 52779 43299
rect 53021 43265 53055 43299
rect 37289 43197 37323 43231
rect 39865 43197 39899 43231
rect 40328 43215 40362 43249
rect 40601 43197 40635 43231
rect 45569 43197 45603 43231
rect 46489 43197 46523 43231
rect 49341 43197 49375 43231
rect 49614 43215 49648 43249
rect 50077 43197 50111 43231
rect 52929 43197 52963 43231
rect 2605 43061 2639 43095
rect 38669 43061 38703 43095
rect 44281 43061 44315 43095
rect 46305 43061 46339 43095
rect 48237 43061 48271 43095
rect 52745 43061 52779 43095
rect 38025 42857 38059 42891
rect 40049 42857 40083 42891
rect 45385 42857 45419 42891
rect 49617 42857 49651 42891
rect 44465 42789 44499 42823
rect 41383 42721 41417 42755
rect 41889 42721 41923 42755
rect 45293 42721 45327 42755
rect 46048 42721 46082 42755
rect 48240 42721 48274 42755
rect 50353 42721 50387 42755
rect 51825 42721 51859 42755
rect 52331 42721 52365 42755
rect 3985 42653 4019 42687
rect 36645 42653 36679 42687
rect 36912 42653 36946 42687
rect 41153 42653 41187 42687
rect 43085 42653 43119 42687
rect 45385 42653 45419 42687
rect 45845 42653 45879 42687
rect 45937 42653 45971 42687
rect 47777 42653 47811 42687
rect 48100 42653 48134 42687
rect 48513 42653 48547 42687
rect 50629 42653 50663 42687
rect 52561 42653 52595 42687
rect 57253 42653 57287 42687
rect 43352 42585 43386 42619
rect 46121 42585 46155 42619
rect 3893 42517 3927 42551
rect 41422 42517 41456 42551
rect 45017 42517 45051 42551
rect 51365 42517 51399 42551
rect 52291 42517 52325 42551
rect 53665 42517 53699 42551
rect 44189 42313 44223 42347
rect 46949 42313 46983 42347
rect 48421 42313 48455 42347
rect 49794 42313 49828 42347
rect 52101 42313 52135 42347
rect 53757 42313 53791 42347
rect 3985 42245 4019 42279
rect 44005 42245 44039 42279
rect 44833 42245 44867 42279
rect 45017 42245 45051 42279
rect 4169 42177 4203 42211
rect 44281 42177 44315 42211
rect 45109 42177 45143 42211
rect 45825 42177 45859 42211
rect 51365 42177 51399 42211
rect 53021 42177 53055 42211
rect 56885 42177 56919 42211
rect 2789 42109 2823 42143
rect 45569 42109 45603 42143
rect 49525 42109 49559 42143
rect 49798 42109 49832 42143
rect 50261 42109 50295 42143
rect 51089 42109 51123 42143
rect 52745 42109 52779 42143
rect 44005 42041 44039 42075
rect 44833 42041 44867 42075
rect 56793 41973 56827 42007
rect 45109 41769 45143 41803
rect 47133 41769 47167 41803
rect 52745 41769 52779 41803
rect 45753 41633 45787 41667
rect 51733 41633 51767 41667
rect 56333 41633 56367 41667
rect 56517 41633 56551 41667
rect 58173 41633 58207 41667
rect 45017 41565 45051 41599
rect 45201 41565 45235 41599
rect 46020 41565 46054 41599
rect 52009 41565 52043 41599
rect 45753 41225 45787 41259
rect 45569 41089 45603 41123
rect 45753 41089 45787 41123
rect 2421 35037 2455 35071
rect 3985 35037 4019 35071
rect 3893 34901 3927 34935
rect 2145 34629 2179 34663
rect 3801 34629 3835 34663
rect 3985 34493 4019 34527
rect 57069 31841 57103 31875
rect 58173 31773 58207 31807
rect 56977 29121 57011 29155
rect 57069 28985 57103 29019
rect 58081 28917 58115 28951
rect 57713 28577 57747 28611
rect 57989 28577 58023 28611
rect 58173 28577 58207 28611
rect 8217 25993 8251 26027
rect 8309 25857 8343 25891
rect 8953 24769 8987 24803
rect 55597 24769 55631 24803
rect 57069 24769 57103 24803
rect 9965 24701 9999 24735
rect 56241 24701 56275 24735
rect 56977 24565 57011 24599
rect 57897 24565 57931 24599
rect 56333 24225 56367 24259
rect 56517 24225 56551 24259
rect 58173 24225 58207 24259
rect 57069 23749 57103 23783
rect 55597 23477 55631 23511
rect 8217 23137 8251 23171
rect 7757 23069 7791 23103
rect 7573 22593 7607 22627
rect 8861 22389 8895 22423
rect 56333 19329 56367 19363
rect 56425 19125 56459 19159
rect 57897 19125 57931 19159
rect 56333 18785 56367 18819
rect 56517 18785 56551 18819
rect 58173 18785 58207 18819
rect 57253 12189 57287 12223
rect 56977 11713 57011 11747
rect 57069 11509 57103 11543
rect 56333 11169 56367 11203
rect 56517 11169 56551 11203
rect 58173 11169 58207 11203
rect 2513 11101 2547 11135
rect 2421 10965 2455 10999
rect 2145 10693 2179 10727
rect 1961 10557 1995 10591
rect 2789 10557 2823 10591
rect 2053 10217 2087 10251
rect 56333 8993 56367 9027
rect 56517 8857 56551 8891
rect 58173 8857 58207 8891
rect 56425 8585 56459 8619
rect 56333 8449 56367 8483
rect 57897 8449 57931 8483
rect 2053 4981 2087 5015
rect 2513 4573 2547 4607
rect 56333 4573 56367 4607
rect 56517 4505 56551 4539
rect 58173 4505 58207 4539
rect 2421 4437 2455 4471
rect 2145 4165 2179 4199
rect 1961 4097 1995 4131
rect 7573 4097 7607 4131
rect 57897 4097 57931 4131
rect 2789 4029 2823 4063
rect 8769 4029 8803 4063
rect 56885 4029 56919 4063
rect 57161 4029 57195 4063
rect 57345 4029 57379 4063
rect 57989 3961 58023 3995
rect 4261 3893 4295 3927
rect 20729 3893 20763 3927
rect 51549 3893 51583 3927
rect 54493 3893 54527 3927
rect 55781 3689 55815 3723
rect 4077 3553 4111 3587
rect 4629 3553 4663 3587
rect 14933 3553 14967 3587
rect 45477 3553 45511 3587
rect 51549 3553 51583 3587
rect 52193 3553 52227 3587
rect 57897 3553 57931 3587
rect 7573 3485 7607 3519
rect 14473 3485 14507 3519
rect 18705 3485 18739 3519
rect 20637 3485 20671 3519
rect 44281 3485 44315 3519
rect 45017 3485 45051 3519
rect 54585 3485 54619 3519
rect 55689 3485 55723 3519
rect 56333 3485 56367 3519
rect 4261 3417 4295 3451
rect 8217 3417 8251 3451
rect 14657 3417 14691 3451
rect 16865 3417 16899 3451
rect 18521 3417 18555 3451
rect 20821 3417 20855 3451
rect 22477 3417 22511 3451
rect 44373 3417 44407 3451
rect 45201 3417 45235 3451
rect 51733 3417 51767 3451
rect 56517 3417 56551 3451
rect 54677 3349 54711 3383
rect 4261 3145 4295 3179
rect 15485 3145 15519 3179
rect 18429 3145 18463 3179
rect 20821 3145 20855 3179
rect 51641 3145 51675 3179
rect 56885 3145 56919 3179
rect 54677 3077 54711 3111
rect 4169 3009 4203 3043
rect 14473 3009 14507 3043
rect 15577 3009 15611 3043
rect 17417 3009 17451 3043
rect 18521 3009 18555 3043
rect 20729 3009 20763 3043
rect 44649 3009 44683 3043
rect 51549 3009 51583 3043
rect 54493 3009 54527 3043
rect 56793 3009 56827 3043
rect 57897 3009 57931 3043
rect 54953 2941 54987 2975
rect 7573 2601 7607 2635
rect 56793 2601 56827 2635
rect 57897 2533 57931 2567
rect 24501 2397 24535 2431
rect 7297 2329 7331 2363
rect 25053 2329 25087 2363
<< metal1 >>
rect 1104 57690 58880 57712
rect 1104 57638 19574 57690
rect 19626 57638 19638 57690
rect 19690 57638 19702 57690
rect 19754 57638 19766 57690
rect 19818 57638 19830 57690
rect 19882 57638 50294 57690
rect 50346 57638 50358 57690
rect 50410 57638 50422 57690
rect 50474 57638 50486 57690
rect 50538 57638 50550 57690
rect 50602 57638 58880 57690
rect 1104 57616 58880 57638
rect 41049 57443 41107 57449
rect 41049 57409 41061 57443
rect 41095 57440 41107 57443
rect 41230 57440 41236 57452
rect 41095 57412 41236 57440
rect 41095 57409 41107 57412
rect 41049 57403 41107 57409
rect 41230 57400 41236 57412
rect 41288 57400 41294 57452
rect 41690 57372 41696 57384
rect 41651 57344 41696 57372
rect 41690 57332 41696 57344
rect 41748 57332 41754 57384
rect 1104 57146 58880 57168
rect 1104 57094 4214 57146
rect 4266 57094 4278 57146
rect 4330 57094 4342 57146
rect 4394 57094 4406 57146
rect 4458 57094 4470 57146
rect 4522 57094 34934 57146
rect 34986 57094 34998 57146
rect 35050 57094 35062 57146
rect 35114 57094 35126 57146
rect 35178 57094 35190 57146
rect 35242 57094 58880 57146
rect 1104 57072 58880 57094
rect 7837 56831 7895 56837
rect 7837 56797 7849 56831
rect 7883 56828 7895 56831
rect 8478 56828 8484 56840
rect 7883 56800 8484 56828
rect 7883 56797 7895 56800
rect 7837 56791 7895 56797
rect 8478 56788 8484 56800
rect 8536 56788 8542 56840
rect 8938 56788 8944 56840
rect 8996 56828 9002 56840
rect 9033 56831 9091 56837
rect 9033 56828 9045 56831
rect 8996 56800 9045 56828
rect 8996 56788 9002 56800
rect 9033 56797 9045 56800
rect 9079 56797 9091 56831
rect 9033 56791 9091 56797
rect 25958 56788 25964 56840
rect 26016 56828 26022 56840
rect 26053 56831 26111 56837
rect 26053 56828 26065 56831
rect 26016 56800 26065 56828
rect 26016 56788 26022 56800
rect 26053 56797 26065 56800
rect 26099 56797 26111 56831
rect 26053 56791 26111 56797
rect 33502 56788 33508 56840
rect 33560 56828 33566 56840
rect 33597 56831 33655 56837
rect 33597 56828 33609 56831
rect 33560 56800 33609 56828
rect 33560 56788 33566 56800
rect 33597 56797 33609 56800
rect 33643 56797 33655 56831
rect 35710 56828 35716 56840
rect 35671 56800 35716 56828
rect 33597 56791 33655 56797
rect 35710 56788 35716 56800
rect 35768 56788 35774 56840
rect 42518 56828 42524 56840
rect 42479 56800 42524 56828
rect 42518 56788 42524 56800
rect 42576 56788 42582 56840
rect 43162 56828 43168 56840
rect 43123 56800 43168 56828
rect 43162 56788 43168 56800
rect 43220 56788 43226 56840
rect 49878 56788 49884 56840
rect 49936 56828 49942 56840
rect 50157 56831 50215 56837
rect 50157 56828 50169 56831
rect 49936 56800 50169 56828
rect 49936 56788 49942 56800
rect 50157 56797 50169 56800
rect 50203 56797 50215 56831
rect 50157 56791 50215 56797
rect 52822 56788 52828 56840
rect 52880 56828 52886 56840
rect 52917 56831 52975 56837
rect 52917 56828 52929 56831
rect 52880 56800 52929 56828
rect 52880 56788 52886 56800
rect 52917 56797 52929 56800
rect 52963 56797 52975 56831
rect 52917 56791 52975 56797
rect 1104 56602 58880 56624
rect 1104 56550 19574 56602
rect 19626 56550 19638 56602
rect 19690 56550 19702 56602
rect 19754 56550 19766 56602
rect 19818 56550 19830 56602
rect 19882 56550 50294 56602
rect 50346 56550 50358 56602
rect 50410 56550 50422 56602
rect 50474 56550 50486 56602
rect 50538 56550 50550 56602
rect 50602 56550 58880 56602
rect 1104 56528 58880 56550
rect 658 56380 664 56432
rect 716 56420 722 56432
rect 43257 56423 43315 56429
rect 43257 56420 43269 56423
rect 716 56392 43269 56420
rect 716 56380 722 56392
rect 43257 56389 43269 56392
rect 43303 56389 43315 56423
rect 43257 56383 43315 56389
rect 8478 56312 8484 56364
rect 8536 56352 8542 56364
rect 8938 56352 8944 56364
rect 8536 56324 8581 56352
rect 8899 56324 8944 56352
rect 8536 56312 8542 56324
rect 8938 56312 8944 56324
rect 8996 56312 9002 56364
rect 33502 56352 33508 56364
rect 33463 56324 33508 56352
rect 33502 56312 33508 56324
rect 33560 56312 33566 56364
rect 49878 56352 49884 56364
rect 49839 56324 49884 56352
rect 49878 56312 49884 56324
rect 49936 56312 49942 56364
rect 52822 56352 52828 56364
rect 52783 56324 52828 56352
rect 52822 56312 52828 56324
rect 52880 56312 52886 56364
rect 7742 56284 7748 56296
rect 7703 56256 7748 56284
rect 7742 56244 7748 56256
rect 7800 56244 7806 56296
rect 8202 56244 8208 56296
rect 8260 56284 8266 56296
rect 8297 56287 8355 56293
rect 8297 56284 8309 56287
rect 8260 56256 8309 56284
rect 8260 56244 8266 56256
rect 8297 56253 8309 56256
rect 8343 56253 8355 56287
rect 9122 56284 9128 56296
rect 9083 56256 9128 56284
rect 8297 56247 8355 56253
rect 9122 56244 9128 56256
rect 9180 56244 9186 56296
rect 9674 56284 9680 56296
rect 9635 56256 9680 56284
rect 9674 56244 9680 56256
rect 9732 56244 9738 56296
rect 33686 56284 33692 56296
rect 33647 56256 33692 56284
rect 33686 56244 33692 56256
rect 33744 56244 33750 56296
rect 34146 56284 34152 56296
rect 34107 56256 34152 56284
rect 34146 56244 34152 56256
rect 34204 56244 34210 56296
rect 44358 56244 44364 56296
rect 44416 56284 44422 56296
rect 44913 56287 44971 56293
rect 44913 56284 44925 56287
rect 44416 56256 44925 56284
rect 44416 56244 44422 56256
rect 44913 56253 44925 56256
rect 44959 56253 44971 56287
rect 45094 56284 45100 56296
rect 45055 56256 45100 56284
rect 44913 56247 44971 56253
rect 45094 56244 45100 56256
rect 45152 56244 45158 56296
rect 50065 56287 50123 56293
rect 50065 56253 50077 56287
rect 50111 56284 50123 56287
rect 50246 56284 50252 56296
rect 50111 56256 50252 56284
rect 50111 56253 50123 56256
rect 50065 56247 50123 56253
rect 50246 56244 50252 56256
rect 50304 56244 50310 56296
rect 50890 56244 50896 56296
rect 50948 56284 50954 56296
rect 51077 56287 51135 56293
rect 51077 56284 51089 56287
rect 50948 56256 51089 56284
rect 50948 56244 50954 56256
rect 51077 56253 51089 56256
rect 51123 56253 51135 56287
rect 51077 56247 51135 56253
rect 53009 56287 53067 56293
rect 53009 56253 53021 56287
rect 53055 56284 53067 56287
rect 53190 56284 53196 56296
rect 53055 56256 53196 56284
rect 53055 56253 53067 56256
rect 53009 56247 53067 56253
rect 53190 56244 53196 56256
rect 53248 56244 53254 56296
rect 53285 56287 53343 56293
rect 53285 56253 53297 56287
rect 53331 56253 53343 56287
rect 53285 56247 53343 56253
rect 26050 56176 26056 56228
rect 26108 56216 26114 56228
rect 50338 56216 50344 56228
rect 26108 56188 50344 56216
rect 26108 56176 26114 56188
rect 50338 56176 50344 56188
rect 50396 56176 50402 56228
rect 52914 56176 52920 56228
rect 52972 56216 52978 56228
rect 53300 56216 53328 56247
rect 52972 56188 53328 56216
rect 52972 56176 52978 56188
rect 42613 56151 42671 56157
rect 42613 56117 42625 56151
rect 42659 56148 42671 56151
rect 43714 56148 43720 56160
rect 42659 56120 43720 56148
rect 42659 56117 42671 56120
rect 42613 56111 42671 56117
rect 43714 56108 43720 56120
rect 43772 56108 43778 56160
rect 1104 56058 58880 56080
rect 1104 56006 4214 56058
rect 4266 56006 4278 56058
rect 4330 56006 4342 56058
rect 4394 56006 4406 56058
rect 4458 56006 4470 56058
rect 4522 56006 34934 56058
rect 34986 56006 34998 56058
rect 35050 56006 35062 56058
rect 35114 56006 35126 56058
rect 35178 56006 35190 56058
rect 35242 56006 58880 56058
rect 1104 55984 58880 56006
rect 33686 55944 33692 55956
rect 33647 55916 33692 55944
rect 33686 55904 33692 55916
rect 33744 55904 33750 55956
rect 44358 55944 44364 55956
rect 35866 55916 43392 55944
rect 44319 55916 44364 55944
rect 35866 55876 35894 55916
rect 33612 55848 35894 55876
rect 25958 55808 25964 55820
rect 25919 55780 25964 55808
rect 25958 55768 25964 55780
rect 26016 55768 26022 55820
rect 26418 55808 26424 55820
rect 26379 55780 26424 55808
rect 26418 55768 26424 55780
rect 26476 55768 26482 55820
rect 33612 55752 33640 55848
rect 35710 55808 35716 55820
rect 35671 55780 35716 55808
rect 35710 55768 35716 55780
rect 35768 55768 35774 55820
rect 36078 55768 36084 55820
rect 36136 55808 36142 55820
rect 36173 55811 36231 55817
rect 36173 55808 36185 55811
rect 36136 55780 36185 55808
rect 36136 55768 36142 55780
rect 36173 55777 36185 55780
rect 36219 55777 36231 55811
rect 36173 55771 36231 55777
rect 41690 55768 41696 55820
rect 41748 55808 41754 55820
rect 41969 55811 42027 55817
rect 41969 55808 41981 55811
rect 41748 55780 41981 55808
rect 41748 55768 41754 55780
rect 41969 55777 41981 55780
rect 42015 55777 42027 55811
rect 41969 55771 42027 55777
rect 42432 55811 42490 55817
rect 42432 55777 42444 55811
rect 42478 55808 42490 55811
rect 42518 55808 42524 55820
rect 42478 55780 42524 55808
rect 42478 55777 42490 55780
rect 42432 55771 42490 55777
rect 42518 55768 42524 55780
rect 42576 55768 42582 55820
rect 43364 55808 43392 55916
rect 44358 55904 44364 55916
rect 44416 55904 44422 55956
rect 50246 55944 50252 55956
rect 50207 55916 50252 55944
rect 50246 55904 50252 55916
rect 50304 55904 50310 55956
rect 53190 55944 53196 55956
rect 53151 55916 53196 55944
rect 53190 55904 53196 55916
rect 53248 55904 53254 55956
rect 43364 55780 53328 55808
rect 33594 55740 33600 55752
rect 33507 55712 33600 55740
rect 33594 55700 33600 55712
rect 33652 55700 33658 55752
rect 42702 55740 42708 55752
rect 42663 55712 42708 55740
rect 42702 55700 42708 55712
rect 42760 55700 42766 55752
rect 43438 55700 43444 55752
rect 43496 55740 43502 55752
rect 44453 55743 44511 55749
rect 44453 55740 44465 55743
rect 43496 55712 44465 55740
rect 43496 55700 43502 55712
rect 44453 55709 44465 55712
rect 44499 55740 44511 55743
rect 49694 55740 49700 55752
rect 44499 55712 49700 55740
rect 44499 55709 44511 55712
rect 44453 55703 44511 55709
rect 49694 55700 49700 55712
rect 49752 55700 49758 55752
rect 50338 55700 50344 55752
rect 50396 55751 50402 55752
rect 50396 55742 50407 55751
rect 53300 55749 53328 55780
rect 53285 55743 53343 55749
rect 50396 55740 50568 55742
rect 50396 55714 51396 55740
rect 50396 55705 50407 55714
rect 50540 55712 51396 55714
rect 50396 55700 50402 55705
rect 26142 55672 26148 55684
rect 26103 55644 26148 55672
rect 26142 55632 26148 55644
rect 26200 55632 26206 55684
rect 35894 55632 35900 55684
rect 35952 55672 35958 55684
rect 51368 55672 51396 55712
rect 53285 55709 53297 55743
rect 53331 55740 53343 55743
rect 56870 55740 56876 55752
rect 53331 55712 56876 55740
rect 53331 55709 53343 55712
rect 53285 55703 53343 55709
rect 56870 55700 56876 55712
rect 56928 55700 56934 55752
rect 55582 55672 55588 55684
rect 35952 55644 35997 55672
rect 51368 55644 55588 55672
rect 35952 55632 35958 55644
rect 55582 55632 55588 55644
rect 55640 55632 55646 55684
rect 42435 55607 42493 55613
rect 42435 55573 42447 55607
rect 42481 55604 42493 55607
rect 42978 55604 42984 55616
rect 42481 55576 42984 55604
rect 42481 55573 42493 55576
rect 42435 55567 42493 55573
rect 42978 55564 42984 55576
rect 43036 55564 43042 55616
rect 43070 55564 43076 55616
rect 43128 55604 43134 55616
rect 43809 55607 43867 55613
rect 43809 55604 43821 55607
rect 43128 55576 43821 55604
rect 43128 55564 43134 55576
rect 43809 55573 43821 55576
rect 43855 55573 43867 55607
rect 43809 55567 43867 55573
rect 1104 55514 58880 55536
rect 1104 55462 19574 55514
rect 19626 55462 19638 55514
rect 19690 55462 19702 55514
rect 19754 55462 19766 55514
rect 19818 55462 19830 55514
rect 19882 55462 50294 55514
rect 50346 55462 50358 55514
rect 50410 55462 50422 55514
rect 50474 55462 50486 55514
rect 50538 55462 50550 55514
rect 50602 55462 58880 55514
rect 1104 55440 58880 55462
rect 9122 55400 9128 55412
rect 9083 55372 9128 55400
rect 9122 55360 9128 55372
rect 9180 55360 9186 55412
rect 26142 55400 26148 55412
rect 26103 55372 26148 55400
rect 26142 55360 26148 55372
rect 26200 55360 26206 55412
rect 35894 55360 35900 55412
rect 35952 55400 35958 55412
rect 42429 55403 42487 55409
rect 35952 55372 35997 55400
rect 35952 55360 35958 55372
rect 42429 55369 42441 55403
rect 42475 55400 42487 55403
rect 42702 55400 42708 55412
rect 42475 55372 42708 55400
rect 42475 55369 42487 55372
rect 42429 55363 42487 55369
rect 42702 55360 42708 55372
rect 42760 55360 42766 55412
rect 43530 55360 43536 55412
rect 43588 55400 43594 55412
rect 43802 55403 43860 55409
rect 43802 55400 43814 55403
rect 43588 55372 43814 55400
rect 43588 55360 43594 55372
rect 43802 55369 43814 55372
rect 43848 55369 43860 55403
rect 43802 55363 43860 55369
rect 49694 55360 49700 55412
rect 49752 55400 49758 55412
rect 56226 55400 56232 55412
rect 49752 55372 56232 55400
rect 49752 55360 49758 55372
rect 56226 55360 56232 55372
rect 56284 55360 56290 55412
rect 9030 55264 9036 55276
rect 8991 55236 9036 55264
rect 9030 55224 9036 55236
rect 9088 55224 9094 55276
rect 26050 55264 26056 55276
rect 26011 55236 26056 55264
rect 26050 55224 26056 55236
rect 26108 55224 26114 55276
rect 35805 55267 35863 55273
rect 35805 55233 35817 55267
rect 35851 55264 35863 55267
rect 43438 55264 43444 55276
rect 35851 55236 43444 55264
rect 35851 55233 35863 55236
rect 35805 55227 35863 55233
rect 43438 55224 43444 55236
rect 43496 55224 43502 55276
rect 43533 55267 43591 55273
rect 43533 55233 43545 55267
rect 43579 55264 43591 55267
rect 44174 55264 44180 55276
rect 43579 55236 44180 55264
rect 43579 55233 43591 55236
rect 43533 55227 43591 55233
rect 44174 55224 44180 55236
rect 44232 55224 44238 55276
rect 44269 55267 44327 55273
rect 44269 55233 44281 55267
rect 44315 55233 44327 55267
rect 44269 55227 44327 55233
rect 43714 55156 43720 55208
rect 43772 55196 43778 55208
rect 43806 55199 43864 55205
rect 43806 55196 43818 55199
rect 43772 55168 43818 55196
rect 43772 55156 43778 55168
rect 43806 55165 43818 55168
rect 43852 55165 43864 55199
rect 43806 55159 43864 55165
rect 42334 55020 42340 55072
rect 42392 55060 42398 55072
rect 44284 55060 44312 55227
rect 42392 55032 44312 55060
rect 42392 55020 42398 55032
rect 1104 54970 58880 54992
rect 1104 54918 4214 54970
rect 4266 54918 4278 54970
rect 4330 54918 4342 54970
rect 4394 54918 4406 54970
rect 4458 54918 4470 54970
rect 4522 54918 34934 54970
rect 34986 54918 34998 54970
rect 35050 54918 35062 54970
rect 35114 54918 35126 54970
rect 35178 54918 35190 54970
rect 35242 54918 58880 54970
rect 1104 54896 58880 54918
rect 44177 54859 44235 54865
rect 44177 54825 44189 54859
rect 44223 54856 44235 54859
rect 45094 54856 45100 54868
rect 44223 54828 45100 54856
rect 44223 54825 44235 54828
rect 44177 54819 44235 54825
rect 45094 54816 45100 54828
rect 45152 54816 45158 54868
rect 41690 54680 41696 54732
rect 41748 54720 41754 54732
rect 42334 54720 42340 54732
rect 41748 54692 42340 54720
rect 41748 54680 41754 54692
rect 42334 54680 42340 54692
rect 42392 54680 42398 54732
rect 42843 54723 42901 54729
rect 42843 54689 42855 54723
rect 42889 54720 42901 54723
rect 43162 54720 43168 54732
rect 42889 54692 43168 54720
rect 42889 54689 42901 54692
rect 42843 54683 42901 54689
rect 43162 54680 43168 54692
rect 43220 54680 43226 54732
rect 1946 54612 1952 54664
rect 2004 54652 2010 54664
rect 2041 54655 2099 54661
rect 2041 54652 2053 54655
rect 2004 54624 2053 54652
rect 2004 54612 2010 54624
rect 2041 54621 2053 54624
rect 2087 54621 2099 54655
rect 43070 54652 43076 54664
rect 43031 54624 43076 54652
rect 2041 54615 2099 54621
rect 43070 54612 43076 54624
rect 43128 54612 43134 54664
rect 42803 54519 42861 54525
rect 42803 54485 42815 54519
rect 42849 54516 42861 54519
rect 42978 54516 42984 54528
rect 42849 54488 42984 54516
rect 42849 54485 42861 54488
rect 42803 54479 42861 54485
rect 42978 54476 42984 54488
rect 43036 54516 43042 54528
rect 43530 54516 43536 54528
rect 43036 54488 43536 54516
rect 43036 54476 43042 54488
rect 43530 54476 43536 54488
rect 43588 54476 43594 54528
rect 1104 54426 58880 54448
rect 1104 54374 19574 54426
rect 19626 54374 19638 54426
rect 19690 54374 19702 54426
rect 19754 54374 19766 54426
rect 19818 54374 19830 54426
rect 19882 54374 50294 54426
rect 50346 54374 50358 54426
rect 50410 54374 50422 54426
rect 50474 54374 50486 54426
rect 50538 54374 50550 54426
rect 50602 54374 58880 54426
rect 1104 54352 58880 54374
rect 1946 54176 1952 54188
rect 1907 54148 1952 54176
rect 1946 54136 1952 54148
rect 2004 54136 2010 54188
rect 46293 54179 46351 54185
rect 46293 54145 46305 54179
rect 46339 54145 46351 54179
rect 46474 54176 46480 54188
rect 46435 54148 46480 54176
rect 46293 54139 46351 54145
rect 2130 54108 2136 54120
rect 2091 54080 2136 54108
rect 2130 54068 2136 54080
rect 2188 54068 2194 54120
rect 2774 54108 2780 54120
rect 2735 54080 2780 54108
rect 2774 54068 2780 54080
rect 2832 54068 2838 54120
rect 46308 54108 46336 54139
rect 46474 54136 46480 54148
rect 46532 54136 46538 54188
rect 47670 54108 47676 54120
rect 46308 54080 47676 54108
rect 47670 54068 47676 54080
rect 47728 54068 47734 54120
rect 46290 53972 46296 53984
rect 46251 53944 46296 53972
rect 46290 53932 46296 53944
rect 46348 53932 46354 53984
rect 1104 53882 58880 53904
rect 1104 53830 4214 53882
rect 4266 53830 4278 53882
rect 4330 53830 4342 53882
rect 4394 53830 4406 53882
rect 4458 53830 4470 53882
rect 4522 53830 34934 53882
rect 34986 53830 34998 53882
rect 35050 53830 35062 53882
rect 35114 53830 35126 53882
rect 35178 53830 35190 53882
rect 35242 53830 58880 53882
rect 1104 53808 58880 53830
rect 2130 53728 2136 53780
rect 2188 53768 2194 53780
rect 2409 53771 2467 53777
rect 2409 53768 2421 53771
rect 2188 53740 2421 53768
rect 2188 53728 2194 53740
rect 2409 53737 2421 53740
rect 2455 53737 2467 53771
rect 2409 53731 2467 53737
rect 46474 53728 46480 53780
rect 46532 53768 46538 53780
rect 46753 53771 46811 53777
rect 46753 53768 46765 53771
rect 46532 53740 46765 53768
rect 46532 53728 46538 53740
rect 46753 53737 46765 53740
rect 46799 53768 46811 53771
rect 49602 53768 49608 53780
rect 46799 53740 49608 53768
rect 46799 53737 46811 53740
rect 46753 53731 46811 53737
rect 49602 53728 49608 53740
rect 49660 53728 49666 53780
rect 45278 53660 45284 53712
rect 45336 53700 45342 53712
rect 45465 53703 45523 53709
rect 45465 53700 45477 53703
rect 45336 53672 45477 53700
rect 45336 53660 45342 53672
rect 45465 53669 45477 53672
rect 45511 53669 45523 53703
rect 45465 53663 45523 53669
rect 2501 53567 2559 53573
rect 2501 53533 2513 53567
rect 2547 53564 2559 53567
rect 2590 53564 2596 53576
rect 2547 53536 2596 53564
rect 2547 53533 2559 53536
rect 2501 53527 2559 53533
rect 2590 53524 2596 53536
rect 2648 53524 2654 53576
rect 42613 53567 42671 53573
rect 42613 53533 42625 53567
rect 42659 53564 42671 53567
rect 42886 53564 42892 53576
rect 42659 53536 42892 53564
rect 42659 53533 42671 53536
rect 42613 53527 42671 53533
rect 42886 53524 42892 53536
rect 42944 53524 42950 53576
rect 45738 53564 45744 53576
rect 45699 53536 45744 53564
rect 45738 53524 45744 53536
rect 45796 53524 45802 53576
rect 45922 53524 45928 53576
rect 45980 53564 45986 53576
rect 46569 53567 46627 53573
rect 46569 53564 46581 53567
rect 45980 53536 46581 53564
rect 45980 53524 45986 53536
rect 46569 53533 46581 53536
rect 46615 53533 46627 53567
rect 46569 53527 46627 53533
rect 45465 53499 45523 53505
rect 45465 53465 45477 53499
rect 45511 53496 45523 53499
rect 47670 53496 47676 53508
rect 45511 53468 47676 53496
rect 45511 53465 45523 53468
rect 45465 53459 45523 53465
rect 47670 53456 47676 53468
rect 47728 53456 47734 53508
rect 45646 53428 45652 53440
rect 45607 53400 45652 53428
rect 45646 53388 45652 53400
rect 45704 53388 45710 53440
rect 1104 53338 58880 53360
rect 1104 53286 19574 53338
rect 19626 53286 19638 53338
rect 19690 53286 19702 53338
rect 19754 53286 19766 53338
rect 19818 53286 19830 53338
rect 19882 53286 50294 53338
rect 50346 53286 50358 53338
rect 50410 53286 50422 53338
rect 50474 53286 50486 53338
rect 50538 53286 50550 53338
rect 50602 53286 58880 53338
rect 1104 53264 58880 53286
rect 44174 53184 44180 53236
rect 44232 53224 44238 53236
rect 44269 53227 44327 53233
rect 44269 53224 44281 53227
rect 44232 53196 44281 53224
rect 44232 53184 44238 53196
rect 44269 53193 44281 53196
rect 44315 53193 44327 53227
rect 44269 53187 44327 53193
rect 46290 53116 46296 53168
rect 46348 53156 46354 53168
rect 46578 53159 46636 53165
rect 46578 53156 46590 53159
rect 46348 53128 46590 53156
rect 46348 53116 46354 53128
rect 46578 53125 46590 53128
rect 46624 53125 46636 53159
rect 46578 53119 46636 53125
rect 49789 53159 49847 53165
rect 49789 53125 49801 53159
rect 49835 53156 49847 53159
rect 49970 53156 49976 53168
rect 49835 53128 49976 53156
rect 49835 53125 49847 53128
rect 49789 53119 49847 53125
rect 49970 53116 49976 53128
rect 50028 53116 50034 53168
rect 42334 53048 42340 53100
rect 42392 53088 42398 53100
rect 42429 53091 42487 53097
rect 42429 53088 42441 53091
rect 42392 53060 42441 53088
rect 42392 53048 42398 53060
rect 42429 53057 42441 53060
rect 42475 53057 42487 53091
rect 42429 53051 42487 53057
rect 42752 53091 42810 53097
rect 42752 53057 42764 53091
rect 42798 53088 42810 53091
rect 42978 53088 42984 53100
rect 42798 53060 42984 53088
rect 42798 53057 42810 53060
rect 42752 53051 42810 53057
rect 42978 53048 42984 53060
rect 43036 53048 43042 53100
rect 48041 53091 48099 53097
rect 48041 53057 48053 53091
rect 48087 53088 48099 53091
rect 48130 53088 48136 53100
rect 48087 53060 48136 53088
rect 48087 53057 48099 53060
rect 48041 53051 48099 53057
rect 48130 53048 48136 53060
rect 48188 53048 48194 53100
rect 48866 53048 48872 53100
rect 48924 53088 48930 53100
rect 49053 53091 49111 53097
rect 49053 53088 49065 53091
rect 48924 53060 49065 53088
rect 48924 53048 48930 53060
rect 49053 53057 49065 53060
rect 49099 53057 49111 53091
rect 49053 53051 49111 53057
rect 42886 52980 42892 53032
rect 42944 53020 42950 53032
rect 43165 53023 43223 53029
rect 42944 52992 42989 53020
rect 42944 52980 42950 52992
rect 43165 52989 43177 53023
rect 43211 53020 43223 53023
rect 43622 53020 43628 53032
rect 43211 52992 43628 53020
rect 43211 52989 43223 52992
rect 43165 52983 43223 52989
rect 43622 52980 43628 52992
rect 43680 52980 43686 53032
rect 46845 53023 46903 53029
rect 46845 52989 46857 53023
rect 46891 53020 46903 53023
rect 46934 53020 46940 53032
rect 46891 52992 46940 53020
rect 46891 52989 46903 52992
rect 46845 52983 46903 52989
rect 46934 52980 46940 52992
rect 46992 53020 46998 53032
rect 47578 53020 47584 53032
rect 46992 52992 47584 53020
rect 46992 52980 46998 52992
rect 47578 52980 47584 52992
rect 47636 52980 47642 53032
rect 47670 52980 47676 53032
rect 47728 53020 47734 53032
rect 47765 53023 47823 53029
rect 47765 53020 47777 53023
rect 47728 52992 47777 53020
rect 47728 52980 47734 52992
rect 47765 52989 47777 52992
rect 47811 52989 47823 53023
rect 47765 52983 47823 52989
rect 50249 53023 50307 53029
rect 50249 52989 50261 53023
rect 50295 52989 50307 53023
rect 50249 52983 50307 52989
rect 47946 52952 47952 52964
rect 47907 52924 47952 52952
rect 47946 52912 47952 52924
rect 48004 52912 48010 52964
rect 49602 52912 49608 52964
rect 49660 52952 49666 52964
rect 49789 52955 49847 52961
rect 49789 52952 49801 52955
rect 49660 52924 49801 52952
rect 49660 52912 49666 52924
rect 49789 52921 49801 52924
rect 49835 52921 49847 52955
rect 49789 52915 49847 52921
rect 45465 52887 45523 52893
rect 45465 52853 45477 52887
rect 45511 52884 45523 52887
rect 45922 52884 45928 52896
rect 45511 52856 45928 52884
rect 45511 52853 45523 52856
rect 45465 52847 45523 52853
rect 45922 52844 45928 52856
rect 45980 52844 45986 52896
rect 47762 52844 47768 52896
rect 47820 52884 47826 52896
rect 47857 52887 47915 52893
rect 47857 52884 47869 52887
rect 47820 52856 47869 52884
rect 47820 52844 47826 52856
rect 47857 52853 47869 52856
rect 47903 52853 47915 52887
rect 49234 52884 49240 52896
rect 49195 52856 49240 52884
rect 47857 52847 47915 52853
rect 49234 52844 49240 52856
rect 49292 52884 49298 52896
rect 50264 52884 50292 52983
rect 50338 52980 50344 53032
rect 50396 53020 50402 53032
rect 50396 52992 50441 53020
rect 50396 52980 50402 52992
rect 50430 52884 50436 52896
rect 49292 52856 50436 52884
rect 49292 52844 49298 52856
rect 50430 52844 50436 52856
rect 50488 52844 50494 52896
rect 50525 52887 50583 52893
rect 50525 52853 50537 52887
rect 50571 52884 50583 52887
rect 51534 52884 51540 52896
rect 50571 52856 51540 52884
rect 50571 52853 50583 52856
rect 50525 52847 50583 52853
rect 51534 52844 51540 52856
rect 51592 52844 51598 52896
rect 1104 52794 58880 52816
rect 1104 52742 4214 52794
rect 4266 52742 4278 52794
rect 4330 52742 4342 52794
rect 4394 52742 4406 52794
rect 4458 52742 4470 52794
rect 4522 52742 34934 52794
rect 34986 52742 34998 52794
rect 35050 52742 35062 52794
rect 35114 52742 35126 52794
rect 35178 52742 35190 52794
rect 35242 52742 58880 52794
rect 1104 52720 58880 52742
rect 41417 52683 41475 52689
rect 41417 52649 41429 52683
rect 41463 52680 41475 52683
rect 42794 52680 42800 52692
rect 41463 52652 42800 52680
rect 41463 52649 41475 52652
rect 41417 52643 41475 52649
rect 42794 52640 42800 52652
rect 42852 52640 42858 52692
rect 43622 52640 43628 52692
rect 43680 52680 43686 52692
rect 43717 52683 43775 52689
rect 43717 52680 43729 52683
rect 43680 52652 43729 52680
rect 43680 52640 43686 52652
rect 43717 52649 43729 52652
rect 43763 52649 43775 52683
rect 46750 52680 46756 52692
rect 43717 52643 43775 52649
rect 45020 52652 46756 52680
rect 41877 52547 41935 52553
rect 41877 52513 41889 52547
rect 41923 52544 41935 52547
rect 42242 52544 42248 52556
rect 41923 52516 42248 52544
rect 41923 52513 41935 52516
rect 41877 52507 41935 52513
rect 42242 52504 42248 52516
rect 42300 52504 42306 52556
rect 45020 52553 45048 52652
rect 46750 52640 46756 52652
rect 46808 52640 46814 52692
rect 46845 52683 46903 52689
rect 46845 52649 46857 52683
rect 46891 52680 46903 52683
rect 46934 52680 46940 52692
rect 46891 52652 46940 52680
rect 46891 52649 46903 52652
rect 46845 52643 46903 52649
rect 46934 52640 46940 52652
rect 46992 52640 46998 52692
rect 48130 52640 48136 52692
rect 48188 52680 48194 52692
rect 49329 52683 49387 52689
rect 49329 52680 49341 52683
rect 48188 52652 49341 52680
rect 48188 52640 48194 52652
rect 49329 52649 49341 52652
rect 49375 52649 49387 52683
rect 49329 52643 49387 52649
rect 46385 52615 46443 52621
rect 46385 52581 46397 52615
rect 46431 52612 46443 52615
rect 48866 52612 48872 52624
rect 46431 52584 46888 52612
rect 48827 52584 48872 52612
rect 46431 52581 46443 52584
rect 46385 52575 46443 52581
rect 42383 52547 42441 52553
rect 42383 52513 42395 52547
rect 42429 52544 42441 52547
rect 44177 52547 44235 52553
rect 44177 52544 44189 52547
rect 42429 52516 44189 52544
rect 42429 52513 42441 52516
rect 42383 52507 42441 52513
rect 44177 52513 44189 52516
rect 44223 52513 44235 52547
rect 44177 52507 44235 52513
rect 45005 52547 45063 52553
rect 45005 52513 45017 52547
rect 45051 52513 45063 52547
rect 45005 52507 45063 52513
rect 46860 52488 46888 52584
rect 48866 52572 48872 52584
rect 48924 52572 48930 52624
rect 50249 52615 50307 52621
rect 50249 52612 50261 52615
rect 49620 52584 50261 52612
rect 49620 52488 49648 52584
rect 50249 52581 50261 52584
rect 50295 52612 50307 52615
rect 50338 52612 50344 52624
rect 50295 52584 50344 52612
rect 50295 52581 50307 52584
rect 50249 52575 50307 52581
rect 50338 52572 50344 52584
rect 50396 52572 50402 52624
rect 50801 52547 50859 52553
rect 50801 52544 50813 52547
rect 49712 52516 50813 52544
rect 42610 52476 42616 52488
rect 42571 52448 42616 52476
rect 42610 52436 42616 52448
rect 42668 52436 42674 52488
rect 45278 52485 45284 52488
rect 45272 52476 45284 52485
rect 45239 52448 45284 52476
rect 45272 52439 45284 52448
rect 45278 52436 45284 52439
rect 45336 52436 45342 52488
rect 46842 52436 46848 52488
rect 46900 52476 46906 52488
rect 47029 52479 47087 52485
rect 47029 52476 47041 52479
rect 46900 52448 47041 52476
rect 46900 52436 46906 52448
rect 47029 52445 47041 52448
rect 47075 52445 47087 52479
rect 47029 52439 47087 52445
rect 47489 52479 47547 52485
rect 47489 52445 47501 52479
rect 47535 52476 47547 52479
rect 47578 52476 47584 52488
rect 47535 52448 47584 52476
rect 47535 52445 47547 52448
rect 47489 52439 47547 52445
rect 47578 52436 47584 52448
rect 47636 52436 47642 52488
rect 47762 52485 47768 52488
rect 47756 52476 47768 52485
rect 47723 52448 47768 52476
rect 47756 52439 47768 52448
rect 47762 52436 47768 52439
rect 47820 52436 47826 52488
rect 49234 52436 49240 52488
rect 49292 52476 49298 52488
rect 49329 52479 49387 52485
rect 49329 52476 49341 52479
rect 49292 52448 49341 52476
rect 49292 52436 49298 52448
rect 49329 52445 49341 52448
rect 49375 52445 49387 52479
rect 49602 52476 49608 52488
rect 49563 52448 49608 52476
rect 49329 52439 49387 52445
rect 49602 52436 49608 52448
rect 49660 52436 49666 52488
rect 49510 52408 49516 52420
rect 49471 52380 49516 52408
rect 49510 52368 49516 52380
rect 49568 52408 49574 52420
rect 49712 52408 49740 52516
rect 50801 52513 50813 52516
rect 50847 52513 50859 52547
rect 50801 52507 50859 52513
rect 50430 52436 50436 52488
rect 50488 52476 50494 52488
rect 50709 52479 50767 52485
rect 50709 52476 50721 52479
rect 50488 52448 50721 52476
rect 50488 52436 50494 52448
rect 50709 52445 50721 52448
rect 50755 52445 50767 52479
rect 50709 52439 50767 52445
rect 49568 52380 49740 52408
rect 49568 52368 49574 52380
rect 49970 52368 49976 52420
rect 50028 52408 50034 52420
rect 50249 52411 50307 52417
rect 50249 52408 50261 52411
rect 50028 52380 50261 52408
rect 50028 52368 50034 52380
rect 50249 52377 50261 52380
rect 50295 52377 50307 52411
rect 50249 52371 50307 52377
rect 42343 52343 42401 52349
rect 42343 52309 42355 52343
rect 42389 52340 42401 52343
rect 42978 52340 42984 52352
rect 42389 52312 42984 52340
rect 42389 52309 42401 52312
rect 42343 52303 42401 52309
rect 42978 52300 42984 52312
rect 43036 52340 43042 52352
rect 43806 52340 43812 52352
rect 43036 52312 43812 52340
rect 43036 52300 43042 52312
rect 43806 52300 43812 52312
rect 43864 52300 43870 52352
rect 50982 52340 50988 52352
rect 50943 52312 50988 52340
rect 50982 52300 50988 52312
rect 51040 52300 51046 52352
rect 1104 52250 58880 52272
rect 1104 52198 19574 52250
rect 19626 52198 19638 52250
rect 19690 52198 19702 52250
rect 19754 52198 19766 52250
rect 19818 52198 19830 52250
rect 19882 52198 50294 52250
rect 50346 52198 50358 52250
rect 50410 52198 50422 52250
rect 50474 52198 50486 52250
rect 50538 52198 50550 52250
rect 50602 52198 58880 52250
rect 1104 52176 58880 52198
rect 42429 52139 42487 52145
rect 42429 52105 42441 52139
rect 42475 52136 42487 52139
rect 42610 52136 42616 52148
rect 42475 52108 42616 52136
rect 42475 52105 42487 52108
rect 42429 52099 42487 52105
rect 42610 52096 42616 52108
rect 42668 52096 42674 52148
rect 43806 52145 43812 52148
rect 43802 52099 43812 52145
rect 43864 52136 43870 52148
rect 45557 52139 45615 52145
rect 43864 52108 43902 52136
rect 43806 52096 43812 52099
rect 43864 52096 43870 52108
rect 45557 52105 45569 52139
rect 45603 52136 45615 52139
rect 45646 52136 45652 52148
rect 45603 52108 45652 52136
rect 45603 52105 45615 52108
rect 45557 52099 45615 52105
rect 45646 52096 45652 52108
rect 45704 52096 45710 52148
rect 45738 52096 45744 52148
rect 45796 52136 45802 52148
rect 46014 52136 46020 52148
rect 45796 52108 46020 52136
rect 45796 52096 45802 52108
rect 46014 52096 46020 52108
rect 46072 52136 46078 52148
rect 46477 52139 46535 52145
rect 46477 52136 46489 52139
rect 46072 52108 46489 52136
rect 46072 52096 46078 52108
rect 46477 52105 46489 52108
rect 46523 52105 46535 52139
rect 47946 52136 47952 52148
rect 47907 52108 47952 52136
rect 46477 52099 46535 52105
rect 47946 52096 47952 52108
rect 48004 52096 48010 52148
rect 49510 52136 49516 52148
rect 49471 52108 49516 52136
rect 49510 52096 49516 52108
rect 49568 52096 49574 52148
rect 47581 52071 47639 52077
rect 47581 52068 47593 52071
rect 46676 52040 47593 52068
rect 46676 52012 46704 52040
rect 47581 52037 47593 52040
rect 47627 52037 47639 52071
rect 47581 52031 47639 52037
rect 47797 52071 47855 52077
rect 47797 52037 47809 52071
rect 47843 52068 47855 52071
rect 48314 52068 48320 52080
rect 47843 52040 48320 52068
rect 47843 52037 47855 52040
rect 47797 52031 47855 52037
rect 48314 52028 48320 52040
rect 48372 52068 48378 52080
rect 48866 52068 48872 52080
rect 48372 52040 48872 52068
rect 48372 52028 48378 52040
rect 48866 52028 48872 52040
rect 48924 52028 48930 52080
rect 49234 52028 49240 52080
rect 49292 52068 49298 52080
rect 49973 52071 50031 52077
rect 49973 52068 49985 52071
rect 49292 52040 49985 52068
rect 49292 52028 49298 52040
rect 49973 52037 49985 52040
rect 50019 52068 50031 52071
rect 50019 52050 51028 52068
rect 50019 52040 51074 52050
rect 50019 52037 50031 52040
rect 49973 52031 50031 52037
rect 51000 52022 51074 52040
rect 51046 52015 51074 52022
rect 42794 51960 42800 52012
rect 42852 52000 42858 52012
rect 42852 51972 43668 52000
rect 42852 51960 42858 51972
rect 43530 51932 43536 51944
rect 43491 51904 43536 51932
rect 43530 51892 43536 51904
rect 43588 51892 43594 51944
rect 43640 51932 43668 51972
rect 45922 51960 45928 52012
rect 45980 52000 45986 52012
rect 46017 52003 46075 52009
rect 46017 52000 46029 52003
rect 45980 51972 46029 52000
rect 45980 51960 45986 51972
rect 46017 51969 46029 51972
rect 46063 52000 46075 52003
rect 46658 52000 46664 52012
rect 46063 51972 46664 52000
rect 46063 51969 46075 51972
rect 46017 51963 46075 51969
rect 46658 51960 46664 51972
rect 46716 51960 46722 52012
rect 46934 52000 46940 52012
rect 46895 51972 46940 52000
rect 46934 51960 46940 51972
rect 46992 52000 46998 52012
rect 49421 52003 49479 52009
rect 49421 52000 49433 52003
rect 46992 51972 49433 52000
rect 46992 51960 46998 51972
rect 49421 51969 49433 51972
rect 49467 52000 49479 52003
rect 49602 52000 49608 52012
rect 49467 51972 49608 52000
rect 49467 51969 49479 51972
rect 49421 51963 49479 51969
rect 49602 51960 49608 51972
rect 49660 51960 49666 52012
rect 51046 52009 51113 52015
rect 51046 51978 51067 52009
rect 51055 51975 51067 51978
rect 51101 51975 51113 52009
rect 51534 52000 51540 52012
rect 51055 51969 51113 51975
rect 51495 51972 51540 52000
rect 51534 51960 51540 51972
rect 51592 51960 51598 52012
rect 43763 51935 43821 51941
rect 43763 51932 43775 51935
rect 43640 51904 43775 51932
rect 43763 51901 43775 51904
rect 43809 51901 43821 51935
rect 43763 51895 43821 51901
rect 44269 51935 44327 51941
rect 44269 51901 44281 51935
rect 44315 51901 44327 51935
rect 44269 51895 44327 51901
rect 42334 51756 42340 51808
rect 42392 51796 42398 51808
rect 44284 51796 44312 51895
rect 46106 51892 46112 51944
rect 46164 51932 46170 51944
rect 50801 51935 50859 51941
rect 50801 51932 50813 51935
rect 46164 51904 46980 51932
rect 46164 51892 46170 51904
rect 46952 51864 46980 51904
rect 49620 51904 50813 51932
rect 49620 51864 49648 51904
rect 50801 51901 50813 51904
rect 50847 51901 50859 51935
rect 50801 51895 50859 51901
rect 49970 51864 49976 51876
rect 45940 51836 46888 51864
rect 46952 51836 49648 51864
rect 49931 51836 49976 51864
rect 45940 51805 45968 51836
rect 46860 51808 46888 51836
rect 49970 51824 49976 51836
rect 50028 51864 50034 51876
rect 50028 51836 50752 51864
rect 50028 51824 50034 51836
rect 42392 51768 44312 51796
rect 45925 51799 45983 51805
rect 42392 51756 42398 51768
rect 45925 51765 45937 51799
rect 45971 51765 45983 51799
rect 46658 51796 46664 51808
rect 46619 51768 46664 51796
rect 45925 51759 45983 51765
rect 46658 51756 46664 51768
rect 46716 51756 46722 51808
rect 46842 51756 46848 51808
rect 46900 51796 46906 51808
rect 47765 51799 47823 51805
rect 47765 51796 47777 51799
rect 46900 51768 47777 51796
rect 46900 51756 46906 51768
rect 47765 51765 47777 51768
rect 47811 51765 47823 51799
rect 47765 51759 47823 51765
rect 49237 51799 49295 51805
rect 49237 51765 49249 51799
rect 49283 51796 49295 51799
rect 49418 51796 49424 51808
rect 49283 51768 49424 51796
rect 49283 51765 49295 51768
rect 49237 51759 49295 51765
rect 49418 51756 49424 51768
rect 49476 51756 49482 51808
rect 50525 51799 50583 51805
rect 50525 51765 50537 51799
rect 50571 51796 50583 51799
rect 50614 51796 50620 51808
rect 50571 51768 50620 51796
rect 50571 51765 50583 51768
rect 50525 51759 50583 51765
rect 50614 51756 50620 51768
rect 50672 51756 50678 51808
rect 50724 51805 50752 51836
rect 50709 51799 50767 51805
rect 50709 51765 50721 51799
rect 50755 51765 50767 51799
rect 50709 51759 50767 51765
rect 51721 51799 51779 51805
rect 51721 51765 51733 51799
rect 51767 51796 51779 51799
rect 52914 51796 52920 51808
rect 51767 51768 52920 51796
rect 51767 51765 51779 51768
rect 51721 51759 51779 51765
rect 52914 51756 52920 51768
rect 52972 51756 52978 51808
rect 1104 51706 58880 51728
rect 1104 51654 4214 51706
rect 4266 51654 4278 51706
rect 4330 51654 4342 51706
rect 4394 51654 4406 51706
rect 4458 51654 4470 51706
rect 4522 51654 34934 51706
rect 34986 51654 34998 51706
rect 35050 51654 35062 51706
rect 35114 51654 35126 51706
rect 35178 51654 35190 51706
rect 35242 51654 58880 51706
rect 1104 51632 58880 51654
rect 46017 51595 46075 51601
rect 46017 51561 46029 51595
rect 46063 51592 46075 51595
rect 46106 51592 46112 51604
rect 46063 51564 46112 51592
rect 46063 51561 46075 51564
rect 46017 51555 46075 51561
rect 46106 51552 46112 51564
rect 46164 51552 46170 51604
rect 45830 51456 45836 51468
rect 45020 51428 45836 51456
rect 44726 51348 44732 51400
rect 44784 51388 44790 51400
rect 45020 51397 45048 51428
rect 45830 51416 45836 51428
rect 45888 51456 45894 51468
rect 47397 51459 47455 51465
rect 47397 51456 47409 51459
rect 45888 51428 47409 51456
rect 45888 51416 45894 51428
rect 47397 51425 47409 51428
rect 47443 51425 47455 51459
rect 47397 51419 47455 51425
rect 45005 51391 45063 51397
rect 45005 51388 45017 51391
rect 44784 51360 45017 51388
rect 44784 51348 44790 51360
rect 45005 51357 45017 51360
rect 45051 51357 45063 51391
rect 45005 51351 45063 51357
rect 45189 51391 45247 51397
rect 45189 51357 45201 51391
rect 45235 51388 45247 51391
rect 45646 51388 45652 51400
rect 45235 51360 45652 51388
rect 45235 51357 45247 51360
rect 45189 51351 45247 51357
rect 45646 51348 45652 51360
rect 45704 51348 45710 51400
rect 45922 51348 45928 51400
rect 45980 51388 45986 51400
rect 46201 51391 46259 51397
rect 46201 51388 46213 51391
rect 45980 51360 46213 51388
rect 45980 51348 45986 51360
rect 46201 51357 46213 51360
rect 46247 51357 46259 51391
rect 46201 51351 46259 51357
rect 46385 51391 46443 51397
rect 46385 51357 46397 51391
rect 46431 51388 46443 51391
rect 46842 51388 46848 51400
rect 46431 51360 46848 51388
rect 46431 51357 46443 51360
rect 46385 51351 46443 51357
rect 46842 51348 46848 51360
rect 46900 51348 46906 51400
rect 47581 51391 47639 51397
rect 47581 51357 47593 51391
rect 47627 51388 47639 51391
rect 48590 51388 48596 51400
rect 47627 51360 48596 51388
rect 47627 51357 47639 51360
rect 47581 51351 47639 51357
rect 48590 51348 48596 51360
rect 48648 51348 48654 51400
rect 50617 51391 50675 51397
rect 50617 51357 50629 51391
rect 50663 51388 50675 51391
rect 50982 51388 50988 51400
rect 50663 51360 50988 51388
rect 50663 51357 50675 51360
rect 50617 51351 50675 51357
rect 50982 51348 50988 51360
rect 51040 51348 51046 51400
rect 47765 51323 47823 51329
rect 47765 51289 47777 51323
rect 47811 51320 47823 51323
rect 48314 51320 48320 51332
rect 47811 51292 48320 51320
rect 47811 51289 47823 51292
rect 47765 51283 47823 51289
rect 48314 51280 48320 51292
rect 48372 51280 48378 51332
rect 45097 51255 45155 51261
rect 45097 51221 45109 51255
rect 45143 51252 45155 51255
rect 45462 51252 45468 51264
rect 45143 51224 45468 51252
rect 45143 51221 45155 51224
rect 45097 51215 45155 51221
rect 45462 51212 45468 51224
rect 45520 51212 45526 51264
rect 50798 51252 50804 51264
rect 50759 51224 50804 51252
rect 50798 51212 50804 51224
rect 50856 51212 50862 51264
rect 1104 51162 58880 51184
rect 1104 51110 19574 51162
rect 19626 51110 19638 51162
rect 19690 51110 19702 51162
rect 19754 51110 19766 51162
rect 19818 51110 19830 51162
rect 19882 51110 50294 51162
rect 50346 51110 50358 51162
rect 50410 51110 50422 51162
rect 50474 51110 50486 51162
rect 50538 51110 50550 51162
rect 50602 51110 58880 51162
rect 1104 51088 58880 51110
rect 48593 51051 48651 51057
rect 48593 51017 48605 51051
rect 48639 51048 48651 51051
rect 49970 51048 49976 51060
rect 48639 51020 49976 51048
rect 48639 51017 48651 51020
rect 48593 51011 48651 51017
rect 49970 51008 49976 51020
rect 50028 51008 50034 51060
rect 46106 50980 46112 50992
rect 44928 50952 46112 50980
rect 44726 50912 44732 50924
rect 44687 50884 44732 50912
rect 44726 50872 44732 50884
rect 44784 50872 44790 50924
rect 44928 50921 44956 50952
rect 46106 50940 46112 50952
rect 46164 50940 46170 50992
rect 44913 50915 44971 50921
rect 44913 50881 44925 50915
rect 44959 50881 44971 50915
rect 45830 50912 45836 50924
rect 45791 50884 45836 50912
rect 44913 50875 44971 50881
rect 45830 50872 45836 50884
rect 45888 50872 45894 50924
rect 46014 50912 46020 50924
rect 45975 50884 46020 50912
rect 46014 50872 46020 50884
rect 46072 50872 46078 50924
rect 48409 50915 48467 50921
rect 48409 50881 48421 50915
rect 48455 50912 48467 50915
rect 48590 50912 48596 50924
rect 48455 50884 48596 50912
rect 48455 50881 48467 50884
rect 48409 50875 48467 50881
rect 48590 50872 48596 50884
rect 48648 50872 48654 50924
rect 49418 50912 49424 50924
rect 49379 50884 49424 50912
rect 49418 50872 49424 50884
rect 49476 50872 49482 50924
rect 50433 50915 50491 50921
rect 50433 50881 50445 50915
rect 50479 50912 50491 50915
rect 50614 50912 50620 50924
rect 50479 50884 50620 50912
rect 50479 50881 50491 50884
rect 50433 50875 50491 50881
rect 50614 50872 50620 50884
rect 50672 50872 50678 50924
rect 43806 50668 43812 50720
rect 43864 50708 43870 50720
rect 44729 50711 44787 50717
rect 44729 50708 44741 50711
rect 43864 50680 44741 50708
rect 43864 50668 43870 50680
rect 44729 50677 44741 50680
rect 44775 50677 44787 50711
rect 46014 50708 46020 50720
rect 45975 50680 46020 50708
rect 44729 50671 44787 50677
rect 46014 50668 46020 50680
rect 46072 50668 46078 50720
rect 49234 50708 49240 50720
rect 49195 50680 49240 50708
rect 49234 50668 49240 50680
rect 49292 50668 49298 50720
rect 50341 50711 50399 50717
rect 50341 50677 50353 50711
rect 50387 50708 50399 50711
rect 50614 50708 50620 50720
rect 50387 50680 50620 50708
rect 50387 50677 50399 50680
rect 50341 50671 50399 50677
rect 50614 50668 50620 50680
rect 50672 50668 50678 50720
rect 1104 50618 58880 50640
rect 1104 50566 4214 50618
rect 4266 50566 4278 50618
rect 4330 50566 4342 50618
rect 4394 50566 4406 50618
rect 4458 50566 4470 50618
rect 4522 50566 34934 50618
rect 34986 50566 34998 50618
rect 35050 50566 35062 50618
rect 35114 50566 35126 50618
rect 35178 50566 35190 50618
rect 35242 50566 58880 50618
rect 1104 50544 58880 50566
rect 48777 50439 48835 50445
rect 48777 50405 48789 50439
rect 48823 50436 48835 50439
rect 49970 50436 49976 50448
rect 48823 50408 49976 50436
rect 48823 50405 48835 50408
rect 48777 50399 48835 50405
rect 49970 50396 49976 50408
rect 50028 50396 50034 50448
rect 48593 50371 48651 50377
rect 48593 50368 48605 50371
rect 47964 50340 48605 50368
rect 36262 50260 36268 50312
rect 36320 50300 36326 50312
rect 37553 50303 37611 50309
rect 37553 50300 37565 50303
rect 36320 50272 37565 50300
rect 36320 50260 36326 50272
rect 37553 50269 37565 50272
rect 37599 50300 37611 50303
rect 40494 50300 40500 50312
rect 37599 50272 40500 50300
rect 37599 50269 37611 50272
rect 37553 50263 37611 50269
rect 40494 50260 40500 50272
rect 40552 50260 40558 50312
rect 47670 50300 47676 50312
rect 47631 50272 47676 50300
rect 47670 50260 47676 50272
rect 47728 50260 47734 50312
rect 47964 50309 47992 50340
rect 48593 50337 48605 50340
rect 48639 50337 48651 50371
rect 48593 50331 48651 50337
rect 47949 50303 48007 50309
rect 47949 50269 47961 50303
rect 47995 50269 48007 50303
rect 48130 50300 48136 50312
rect 48091 50272 48136 50300
rect 47949 50263 48007 50269
rect 48130 50260 48136 50272
rect 48188 50260 48194 50312
rect 37820 50235 37878 50241
rect 37820 50201 37832 50235
rect 37866 50232 37878 50235
rect 37918 50232 37924 50244
rect 37866 50204 37924 50232
rect 37866 50201 37878 50204
rect 37820 50195 37878 50201
rect 37918 50192 37924 50204
rect 37976 50192 37982 50244
rect 48038 50192 48044 50244
rect 48096 50232 48102 50244
rect 49053 50235 49111 50241
rect 49053 50232 49065 50235
rect 48096 50204 49065 50232
rect 48096 50192 48102 50204
rect 49053 50201 49065 50204
rect 49099 50201 49111 50235
rect 49053 50195 49111 50201
rect 38933 50167 38991 50173
rect 38933 50133 38945 50167
rect 38979 50164 38991 50167
rect 39482 50164 39488 50176
rect 38979 50136 39488 50164
rect 38979 50133 38991 50136
rect 38933 50127 38991 50133
rect 39482 50124 39488 50136
rect 39540 50124 39546 50176
rect 47486 50164 47492 50176
rect 47447 50136 47492 50164
rect 47486 50124 47492 50136
rect 47544 50124 47550 50176
rect 1104 50074 58880 50096
rect 1104 50022 19574 50074
rect 19626 50022 19638 50074
rect 19690 50022 19702 50074
rect 19754 50022 19766 50074
rect 19818 50022 19830 50074
rect 19882 50022 50294 50074
rect 50346 50022 50358 50074
rect 50410 50022 50422 50074
rect 50474 50022 50486 50074
rect 50538 50022 50550 50074
rect 50602 50022 58880 50074
rect 1104 50000 58880 50022
rect 37918 49960 37924 49972
rect 37879 49932 37924 49960
rect 37918 49920 37924 49932
rect 37976 49920 37982 49972
rect 43714 49920 43720 49972
rect 43772 49969 43778 49972
rect 43772 49960 43781 49969
rect 43772 49932 43817 49960
rect 43772 49923 43781 49932
rect 43772 49920 43778 49923
rect 50706 49920 50712 49972
rect 50764 49960 50770 49972
rect 50807 49963 50865 49969
rect 50807 49960 50819 49963
rect 50764 49932 50819 49960
rect 50764 49920 50770 49932
rect 50807 49929 50819 49932
rect 50853 49929 50865 49963
rect 50807 49923 50865 49929
rect 52181 49963 52239 49969
rect 52181 49929 52193 49963
rect 52227 49960 52239 49963
rect 53190 49960 53196 49972
rect 52227 49932 53196 49960
rect 52227 49929 52239 49932
rect 52181 49923 52239 49929
rect 53190 49920 53196 49932
rect 53248 49920 53254 49972
rect 47486 49852 47492 49904
rect 47544 49892 47550 49904
rect 47826 49895 47884 49901
rect 47826 49892 47838 49895
rect 47544 49864 47838 49892
rect 47544 49852 47550 49864
rect 47826 49861 47838 49864
rect 47872 49861 47884 49895
rect 47826 49855 47884 49861
rect 38102 49824 38108 49836
rect 38063 49796 38108 49824
rect 38102 49784 38108 49796
rect 38160 49784 38166 49836
rect 38381 49827 38439 49833
rect 38381 49793 38393 49827
rect 38427 49793 38439 49827
rect 38381 49787 38439 49793
rect 38565 49827 38623 49833
rect 38565 49793 38577 49827
rect 38611 49824 38623 49827
rect 39482 49824 39488 49836
rect 38611 49796 39488 49824
rect 38611 49793 38623 49796
rect 38565 49787 38623 49793
rect 1946 49756 1952 49768
rect 1907 49728 1952 49756
rect 1946 49716 1952 49728
rect 2004 49716 2010 49768
rect 2130 49756 2136 49768
rect 2091 49728 2136 49756
rect 2130 49716 2136 49728
rect 2188 49716 2194 49768
rect 2774 49756 2780 49768
rect 2735 49728 2780 49756
rect 2774 49716 2780 49728
rect 2832 49716 2838 49768
rect 37550 49716 37556 49768
rect 37608 49756 37614 49768
rect 38396 49756 38424 49787
rect 39482 49784 39488 49796
rect 39540 49784 39546 49836
rect 40494 49824 40500 49836
rect 40455 49796 40500 49824
rect 40494 49784 40500 49796
rect 40552 49784 40558 49836
rect 40770 49833 40776 49836
rect 40764 49787 40776 49833
rect 40828 49824 40834 49836
rect 40828 49796 40864 49824
rect 40770 49784 40776 49787
rect 40828 49784 40834 49796
rect 42334 49784 42340 49836
rect 42392 49824 42398 49836
rect 43257 49827 43315 49833
rect 43257 49824 43269 49827
rect 42392 49796 43269 49824
rect 42392 49784 42398 49796
rect 43257 49793 43269 49796
rect 43303 49793 43315 49827
rect 43257 49787 43315 49793
rect 39669 49759 39727 49765
rect 39669 49756 39681 49759
rect 37608 49728 38424 49756
rect 38580 49728 39681 49756
rect 37608 49716 37614 49728
rect 38580 49700 38608 49728
rect 39669 49725 39681 49728
rect 39715 49725 39727 49759
rect 39669 49719 39727 49725
rect 43720 49759 43778 49765
rect 43720 49725 43732 49759
rect 43766 49756 43778 49759
rect 43806 49756 43812 49768
rect 43766 49728 43812 49756
rect 43766 49725 43778 49728
rect 43720 49719 43778 49725
rect 43806 49716 43812 49728
rect 43864 49716 43870 49768
rect 43993 49759 44051 49765
rect 43993 49725 44005 49759
rect 44039 49756 44051 49759
rect 44174 49756 44180 49768
rect 44039 49728 44180 49756
rect 44039 49725 44051 49728
rect 43993 49719 44051 49725
rect 44174 49716 44180 49728
rect 44232 49716 44238 49768
rect 47578 49756 47584 49768
rect 47539 49728 47584 49756
rect 47578 49716 47584 49728
rect 47636 49716 47642 49768
rect 50154 49716 50160 49768
rect 50212 49756 50218 49768
rect 50341 49759 50399 49765
rect 50341 49756 50353 49759
rect 50212 49728 50353 49756
rect 50212 49716 50218 49728
rect 50341 49725 50353 49728
rect 50387 49725 50399 49759
rect 50341 49719 50399 49725
rect 50798 49716 50804 49768
rect 50856 49756 50862 49768
rect 51074 49756 51080 49768
rect 50856 49728 50901 49756
rect 51035 49728 51080 49756
rect 50856 49716 50862 49728
rect 51074 49716 51080 49728
rect 51132 49716 51138 49768
rect 38562 49648 38568 49700
rect 38620 49648 38626 49700
rect 39301 49623 39359 49629
rect 39301 49589 39313 49623
rect 39347 49620 39359 49623
rect 39850 49620 39856 49632
rect 39347 49592 39856 49620
rect 39347 49589 39359 49592
rect 39301 49583 39359 49589
rect 39850 49580 39856 49592
rect 39908 49580 39914 49632
rect 41414 49580 41420 49632
rect 41472 49620 41478 49632
rect 41877 49623 41935 49629
rect 41877 49620 41889 49623
rect 41472 49592 41889 49620
rect 41472 49580 41478 49592
rect 41877 49589 41889 49592
rect 41923 49620 41935 49623
rect 42702 49620 42708 49632
rect 41923 49592 42708 49620
rect 41923 49589 41935 49592
rect 41877 49583 41935 49589
rect 42702 49580 42708 49592
rect 42760 49580 42766 49632
rect 45094 49620 45100 49632
rect 45055 49592 45100 49620
rect 45094 49580 45100 49592
rect 45152 49580 45158 49632
rect 48590 49580 48596 49632
rect 48648 49620 48654 49632
rect 48961 49623 49019 49629
rect 48961 49620 48973 49623
rect 48648 49592 48973 49620
rect 48648 49580 48654 49592
rect 48961 49589 48973 49592
rect 49007 49589 49019 49623
rect 48961 49583 49019 49589
rect 1104 49530 58880 49552
rect 1104 49478 4214 49530
rect 4266 49478 4278 49530
rect 4330 49478 4342 49530
rect 4394 49478 4406 49530
rect 4458 49478 4470 49530
rect 4522 49478 34934 49530
rect 34986 49478 34998 49530
rect 35050 49478 35062 49530
rect 35114 49478 35126 49530
rect 35178 49478 35190 49530
rect 35242 49478 58880 49530
rect 1104 49456 58880 49478
rect 1946 49376 1952 49428
rect 2004 49416 2010 49428
rect 2041 49419 2099 49425
rect 2041 49416 2053 49419
rect 2004 49388 2053 49416
rect 2004 49376 2010 49388
rect 2041 49385 2053 49388
rect 2087 49385 2099 49419
rect 2041 49379 2099 49385
rect 39482 49376 39488 49428
rect 39540 49416 39546 49428
rect 39540 49388 40356 49416
rect 39540 49376 39546 49388
rect 39209 49351 39267 49357
rect 39209 49317 39221 49351
rect 39255 49348 39267 49351
rect 39853 49351 39911 49357
rect 39853 49348 39865 49351
rect 39255 49320 39865 49348
rect 39255 49317 39267 49320
rect 39209 49311 39267 49317
rect 39853 49317 39865 49320
rect 39899 49317 39911 49351
rect 40218 49348 40224 49360
rect 39853 49311 39911 49317
rect 40144 49320 40224 49348
rect 36262 49280 36268 49292
rect 36223 49252 36268 49280
rect 36262 49240 36268 49252
rect 36320 49240 36326 49292
rect 40144 49289 40172 49320
rect 40218 49308 40224 49320
rect 40276 49308 40282 49360
rect 40129 49283 40187 49289
rect 40129 49249 40141 49283
rect 40175 49249 40187 49283
rect 40328 49280 40356 49388
rect 50154 49376 50160 49428
rect 50212 49416 50218 49428
rect 50798 49416 50804 49428
rect 50212 49388 50804 49416
rect 50212 49376 50218 49388
rect 50798 49376 50804 49388
rect 50856 49376 50862 49428
rect 51074 49376 51080 49428
rect 51132 49416 51138 49428
rect 51997 49419 52055 49425
rect 51997 49416 52009 49419
rect 51132 49388 52009 49416
rect 51132 49376 51138 49388
rect 51997 49385 52009 49388
rect 52043 49385 52055 49419
rect 54297 49419 54355 49425
rect 54297 49416 54309 49419
rect 51997 49379 52055 49385
rect 52104 49388 54309 49416
rect 41328 49283 41386 49289
rect 41328 49280 41340 49283
rect 40328 49252 41340 49280
rect 40129 49243 40187 49249
rect 41328 49249 41340 49252
rect 41374 49249 41386 49283
rect 45462 49280 45468 49292
rect 45426 49252 45468 49280
rect 41328 49243 41386 49249
rect 45462 49240 45468 49252
rect 45520 49240 45526 49292
rect 48130 49240 48136 49292
rect 48188 49280 48194 49292
rect 48228 49283 48286 49289
rect 48228 49280 48240 49283
rect 48188 49252 48240 49280
rect 48188 49240 48194 49252
rect 48228 49249 48240 49252
rect 48274 49249 48286 49283
rect 48228 49243 48286 49249
rect 48501 49283 48559 49289
rect 48501 49249 48513 49283
rect 48547 49280 48559 49283
rect 48547 49252 50568 49280
rect 48547 49249 48559 49252
rect 48501 49243 48559 49249
rect 39850 49172 39856 49224
rect 39908 49212 39914 49224
rect 40037 49215 40095 49221
rect 40037 49212 40049 49215
rect 39908 49184 40049 49212
rect 39908 49172 39914 49184
rect 40037 49181 40049 49184
rect 40083 49181 40095 49215
rect 40221 49215 40279 49221
rect 40221 49212 40233 49215
rect 40037 49175 40095 49181
rect 40144 49184 40233 49212
rect 40144 49156 40172 49184
rect 40221 49181 40233 49184
rect 40267 49181 40279 49215
rect 40221 49175 40279 49181
rect 40310 49172 40316 49224
rect 40368 49212 40374 49224
rect 40862 49212 40868 49224
rect 40368 49184 40461 49212
rect 40823 49184 40868 49212
rect 40368 49172 40374 49184
rect 36532 49147 36590 49153
rect 36532 49113 36544 49147
rect 36578 49144 36590 49147
rect 36722 49144 36728 49156
rect 36578 49116 36728 49144
rect 36578 49113 36590 49116
rect 36532 49107 36590 49113
rect 36722 49104 36728 49116
rect 36780 49104 36786 49156
rect 38841 49147 38899 49153
rect 38841 49113 38853 49147
rect 38887 49144 38899 49147
rect 39390 49144 39396 49156
rect 38887 49116 39396 49144
rect 38887 49113 38899 49116
rect 38841 49107 38899 49113
rect 39390 49104 39396 49116
rect 39448 49104 39454 49156
rect 39482 49104 39488 49156
rect 39540 49144 39546 49156
rect 40126 49144 40132 49156
rect 39540 49116 40132 49144
rect 39540 49104 39546 49116
rect 40126 49104 40132 49116
rect 40184 49104 40190 49156
rect 40420 49144 40448 49184
rect 40862 49172 40868 49184
rect 40920 49172 40926 49224
rect 41414 49212 41420 49224
rect 40972 49184 41420 49212
rect 40972 49144 41000 49184
rect 41414 49172 41420 49184
rect 41472 49172 41478 49224
rect 41598 49212 41604 49224
rect 41559 49184 41604 49212
rect 41598 49172 41604 49184
rect 41656 49172 41662 49224
rect 42334 49172 42340 49224
rect 42392 49212 42398 49224
rect 45002 49212 45008 49224
rect 42392 49184 45008 49212
rect 42392 49172 42398 49184
rect 45002 49172 45008 49184
rect 45060 49172 45066 49224
rect 45094 49172 45100 49224
rect 45152 49212 45158 49224
rect 45741 49215 45799 49221
rect 45741 49212 45753 49215
rect 45152 49184 45753 49212
rect 45152 49172 45158 49184
rect 45741 49181 45753 49184
rect 45787 49181 45799 49215
rect 47762 49212 47768 49224
rect 47723 49184 47768 49212
rect 45741 49175 45799 49181
rect 47762 49172 47768 49184
rect 47820 49212 47826 49224
rect 50154 49212 50160 49224
rect 47820 49184 50160 49212
rect 47820 49172 47826 49184
rect 50154 49172 50160 49184
rect 50212 49172 50218 49224
rect 50540 49212 50568 49252
rect 50614 49240 50620 49292
rect 50672 49280 50678 49292
rect 52104 49280 52132 49388
rect 54297 49385 54309 49388
rect 54343 49385 54355 49419
rect 54297 49379 54355 49385
rect 50672 49252 50717 49280
rect 50816 49252 52132 49280
rect 50672 49240 50678 49252
rect 50816 49212 50844 49252
rect 52638 49240 52644 49292
rect 52696 49280 52702 49292
rect 52780 49283 52838 49289
rect 52780 49280 52792 49283
rect 52696 49252 52792 49280
rect 52696 49240 52702 49252
rect 52780 49249 52792 49252
rect 52826 49249 52838 49283
rect 52780 49243 52838 49249
rect 52914 49240 52920 49292
rect 52972 49280 52978 49292
rect 53190 49280 53196 49292
rect 52972 49252 53017 49280
rect 53151 49252 53196 49280
rect 52972 49240 52978 49252
rect 53190 49240 53196 49252
rect 53248 49240 53254 49292
rect 50540 49184 50844 49212
rect 50893 49215 50951 49221
rect 50893 49181 50905 49215
rect 50939 49212 50951 49215
rect 51166 49212 51172 49224
rect 50939 49184 51172 49212
rect 50939 49181 50951 49184
rect 50893 49175 50951 49181
rect 51166 49172 51172 49184
rect 51224 49172 51230 49224
rect 52457 49215 52515 49221
rect 52457 49181 52469 49215
rect 52503 49181 52515 49215
rect 52457 49175 52515 49181
rect 40420 49116 41000 49144
rect 46676 49116 47900 49144
rect 37645 49079 37703 49085
rect 37645 49045 37657 49079
rect 37691 49076 37703 49079
rect 37918 49076 37924 49088
rect 37691 49048 37924 49076
rect 37691 49045 37703 49048
rect 37645 49039 37703 49045
rect 37918 49036 37924 49048
rect 37976 49036 37982 49088
rect 39301 49079 39359 49085
rect 39301 49045 39313 49079
rect 39347 49076 39359 49079
rect 40494 49076 40500 49088
rect 39347 49048 40500 49076
rect 39347 49045 39359 49048
rect 39301 49039 39359 49045
rect 40494 49036 40500 49048
rect 40552 49036 40558 49088
rect 41322 49076 41328 49088
rect 41380 49085 41386 49088
rect 41289 49048 41328 49076
rect 41322 49036 41328 49048
rect 41380 49039 41389 49085
rect 42705 49079 42763 49085
rect 42705 49045 42717 49079
rect 42751 49076 42763 49079
rect 43162 49076 43168 49088
rect 42751 49048 43168 49076
rect 42751 49045 42763 49048
rect 42705 49039 42763 49045
rect 41380 49036 41386 49039
rect 43162 49036 43168 49048
rect 43220 49036 43226 49088
rect 45471 49079 45529 49085
rect 45471 49045 45483 49079
rect 45517 49076 45529 49079
rect 46198 49076 46204 49088
rect 45517 49048 46204 49076
rect 45517 49045 45529 49048
rect 45471 49039 45529 49045
rect 46198 49036 46204 49048
rect 46256 49076 46262 49088
rect 46676 49076 46704 49116
rect 46842 49076 46848 49088
rect 46256 49048 46704 49076
rect 46803 49048 46848 49076
rect 46256 49036 46262 49048
rect 46842 49036 46848 49048
rect 46900 49036 46906 49088
rect 47872 49076 47900 49116
rect 48231 49079 48289 49085
rect 48231 49076 48243 49079
rect 47872 49048 48243 49076
rect 48231 49045 48243 49048
rect 48277 49076 48289 49079
rect 48958 49076 48964 49088
rect 48277 49048 48964 49076
rect 48277 49045 48289 49048
rect 48231 49039 48289 49045
rect 48958 49036 48964 49048
rect 49016 49036 49022 49088
rect 49602 49076 49608 49088
rect 49563 49048 49608 49076
rect 49602 49036 49608 49048
rect 49660 49036 49666 49088
rect 50614 49076 50620 49088
rect 50672 49085 50678 49088
rect 50581 49048 50620 49076
rect 50614 49036 50620 49048
rect 50672 49039 50681 49085
rect 50672 49036 50678 49039
rect 50798 49036 50804 49088
rect 50856 49076 50862 49088
rect 52270 49076 52276 49088
rect 50856 49048 52276 49076
rect 50856 49036 50862 49048
rect 52270 49036 52276 49048
rect 52328 49076 52334 49088
rect 52472 49076 52500 49175
rect 52328 49048 52500 49076
rect 52328 49036 52334 49048
rect 1104 48986 58880 49008
rect 1104 48934 19574 48986
rect 19626 48934 19638 48986
rect 19690 48934 19702 48986
rect 19754 48934 19766 48986
rect 19818 48934 19830 48986
rect 19882 48934 50294 48986
rect 50346 48934 50358 48986
rect 50410 48934 50422 48986
rect 50474 48934 50486 48986
rect 50538 48934 50550 48986
rect 50602 48934 58880 48986
rect 1104 48912 58880 48934
rect 2130 48832 2136 48884
rect 2188 48872 2194 48884
rect 2409 48875 2467 48881
rect 2409 48872 2421 48875
rect 2188 48844 2421 48872
rect 2188 48832 2194 48844
rect 2409 48841 2421 48844
rect 2455 48841 2467 48875
rect 36722 48872 36728 48884
rect 36683 48844 36728 48872
rect 2409 48835 2467 48841
rect 36722 48832 36728 48844
rect 36780 48832 36786 48884
rect 37550 48872 37556 48884
rect 37511 48844 37556 48872
rect 37550 48832 37556 48844
rect 37608 48832 37614 48884
rect 38102 48832 38108 48884
rect 38160 48872 38166 48884
rect 38381 48875 38439 48881
rect 38381 48872 38393 48875
rect 38160 48844 38393 48872
rect 38160 48832 38166 48844
rect 38381 48841 38393 48844
rect 38427 48841 38439 48875
rect 39390 48872 39396 48884
rect 39351 48844 39396 48872
rect 38381 48835 38439 48841
rect 39390 48832 39396 48844
rect 39448 48832 39454 48884
rect 39666 48832 39672 48884
rect 39724 48872 39730 48884
rect 39761 48875 39819 48881
rect 39761 48872 39773 48875
rect 39724 48844 39773 48872
rect 39724 48832 39730 48844
rect 39761 48841 39773 48844
rect 39807 48841 39819 48875
rect 39761 48835 39819 48841
rect 40681 48875 40739 48881
rect 40681 48841 40693 48875
rect 40727 48872 40739 48875
rect 40770 48872 40776 48884
rect 40727 48844 40776 48872
rect 40727 48841 40739 48844
rect 40681 48835 40739 48841
rect 40770 48832 40776 48844
rect 40828 48832 40834 48884
rect 41046 48832 41052 48884
rect 41104 48872 41110 48884
rect 41322 48872 41328 48884
rect 41104 48844 41328 48872
rect 41104 48832 41110 48844
rect 41322 48832 41328 48844
rect 41380 48872 41386 48884
rect 42895 48875 42953 48881
rect 42895 48872 42907 48875
rect 41380 48844 42907 48872
rect 41380 48832 41386 48844
rect 42895 48841 42907 48844
rect 42941 48872 42953 48875
rect 43622 48872 43628 48884
rect 42941 48844 43628 48872
rect 42941 48841 42953 48844
rect 42895 48835 42953 48841
rect 43622 48832 43628 48844
rect 43680 48832 43686 48884
rect 44174 48832 44180 48884
rect 44232 48872 44238 48884
rect 44269 48875 44327 48881
rect 44269 48872 44281 48875
rect 44232 48844 44281 48872
rect 44232 48832 44238 48844
rect 44269 48841 44281 48844
rect 44315 48841 44327 48875
rect 44269 48835 44327 48841
rect 45741 48875 45799 48881
rect 45741 48841 45753 48875
rect 45787 48872 45799 48875
rect 47578 48872 47584 48884
rect 45787 48844 47584 48872
rect 45787 48841 45799 48844
rect 45741 48835 45799 48841
rect 47578 48832 47584 48844
rect 47636 48832 47642 48884
rect 48958 48832 48964 48884
rect 49016 48872 49022 48884
rect 49059 48875 49117 48881
rect 49059 48872 49071 48875
rect 49016 48844 49071 48872
rect 49016 48832 49022 48844
rect 49059 48841 49071 48844
rect 49105 48872 49117 48875
rect 50433 48875 50491 48881
rect 49105 48844 50384 48872
rect 49105 48841 49117 48844
rect 49059 48835 49117 48841
rect 2498 48736 2504 48748
rect 2459 48708 2504 48736
rect 2498 48696 2504 48708
rect 2556 48696 2562 48748
rect 36725 48739 36783 48745
rect 36725 48705 36737 48739
rect 36771 48736 36783 48739
rect 37568 48736 37596 48832
rect 37721 48807 37779 48813
rect 37721 48773 37733 48807
rect 37767 48804 37779 48807
rect 37767 48776 37872 48804
rect 37767 48773 37779 48776
rect 37721 48767 37779 48773
rect 37844 48748 37872 48776
rect 37918 48764 37924 48816
rect 37976 48804 37982 48816
rect 38562 48804 38568 48816
rect 37976 48776 38568 48804
rect 37976 48764 37982 48776
rect 38562 48764 38568 48776
rect 38620 48764 38626 48816
rect 40218 48804 40224 48816
rect 38672 48776 40224 48804
rect 37826 48736 37832 48748
rect 36771 48708 37596 48736
rect 37739 48708 37832 48736
rect 36771 48705 36783 48708
rect 36725 48699 36783 48705
rect 37826 48696 37832 48708
rect 37884 48736 37890 48748
rect 38672 48745 38700 48776
rect 40218 48764 40224 48776
rect 40276 48764 40282 48816
rect 47673 48807 47731 48813
rect 47673 48773 47685 48807
rect 47719 48804 47731 48807
rect 48590 48804 48596 48816
rect 47719 48776 48596 48804
rect 47719 48773 47731 48776
rect 47673 48767 47731 48773
rect 48590 48764 48596 48776
rect 48648 48764 48654 48816
rect 50356 48804 50384 48844
rect 50433 48841 50445 48875
rect 50479 48872 50491 48875
rect 51166 48872 51172 48884
rect 50479 48844 51172 48872
rect 50479 48841 50491 48844
rect 50433 48835 50491 48841
rect 51166 48832 51172 48844
rect 51224 48832 51230 48884
rect 50614 48804 50620 48816
rect 50356 48776 50620 48804
rect 50614 48764 50620 48776
rect 50672 48804 50678 48816
rect 52638 48804 52644 48816
rect 50672 48776 52644 48804
rect 50672 48764 50678 48776
rect 52638 48764 52644 48776
rect 52696 48764 52702 48816
rect 38657 48739 38715 48745
rect 38657 48736 38669 48739
rect 37884 48708 38669 48736
rect 37884 48696 37890 48708
rect 38657 48705 38669 48708
rect 38703 48705 38715 48739
rect 38657 48699 38715 48705
rect 38749 48739 38807 48745
rect 38749 48705 38761 48739
rect 38795 48736 38807 48739
rect 39482 48736 39488 48748
rect 38795 48708 39488 48736
rect 38795 48705 38807 48708
rect 38749 48699 38807 48705
rect 39482 48696 39488 48708
rect 39540 48696 39546 48748
rect 39669 48739 39727 48745
rect 39669 48705 39681 48739
rect 39715 48736 39727 48739
rect 40310 48736 40316 48748
rect 39715 48708 40316 48736
rect 39715 48705 39727 48708
rect 39669 48699 39727 48705
rect 40310 48696 40316 48708
rect 40368 48696 40374 48748
rect 40494 48736 40500 48748
rect 40455 48708 40500 48736
rect 40494 48696 40500 48708
rect 40552 48696 40558 48748
rect 40862 48696 40868 48748
rect 40920 48736 40926 48748
rect 42334 48736 42340 48748
rect 40920 48708 42340 48736
rect 40920 48696 40926 48708
rect 42334 48696 42340 48708
rect 42392 48736 42398 48748
rect 42429 48739 42487 48745
rect 42429 48736 42441 48739
rect 42392 48708 42441 48736
rect 42392 48696 42398 48708
rect 42429 48705 42441 48708
rect 42475 48705 42487 48739
rect 43162 48736 43168 48748
rect 43123 48708 43168 48736
rect 42429 48699 42487 48705
rect 43162 48696 43168 48708
rect 43220 48696 43226 48748
rect 45005 48739 45063 48745
rect 45005 48705 45017 48739
rect 45051 48736 45063 48739
rect 45094 48736 45100 48748
rect 45051 48708 45100 48736
rect 45051 48705 45063 48708
rect 45005 48699 45063 48705
rect 45094 48696 45100 48708
rect 45152 48696 45158 48748
rect 36446 48668 36452 48680
rect 36407 48640 36452 48668
rect 36446 48628 36452 48640
rect 36504 48628 36510 48680
rect 38565 48671 38623 48677
rect 38565 48637 38577 48671
rect 38611 48637 38623 48671
rect 38565 48631 38623 48637
rect 36633 48603 36691 48609
rect 36633 48569 36645 48603
rect 36679 48600 36691 48603
rect 37458 48600 37464 48612
rect 36679 48572 37464 48600
rect 36679 48569 36691 48572
rect 36633 48563 36691 48569
rect 37458 48560 37464 48572
rect 37516 48560 37522 48612
rect 38580 48600 38608 48631
rect 38838 48628 38844 48680
rect 38896 48668 38902 48680
rect 39577 48671 39635 48677
rect 39577 48668 39589 48671
rect 38896 48640 39589 48668
rect 38896 48628 38902 48640
rect 39577 48637 39589 48640
rect 39623 48637 39635 48671
rect 39942 48668 39948 48680
rect 39903 48640 39948 48668
rect 39577 48631 39635 48637
rect 39942 48628 39948 48640
rect 40000 48628 40006 48680
rect 40037 48671 40095 48677
rect 40037 48637 40049 48671
rect 40083 48637 40095 48671
rect 40037 48631 40095 48637
rect 39850 48600 39856 48612
rect 38580 48572 39856 48600
rect 39850 48560 39856 48572
rect 39908 48600 39914 48612
rect 40052 48600 40080 48631
rect 42886 48628 42892 48680
rect 42944 48668 42950 48680
rect 44726 48668 44732 48680
rect 42944 48640 42989 48668
rect 44687 48640 44732 48668
rect 42944 48628 42950 48640
rect 44726 48628 44732 48640
rect 44784 48628 44790 48680
rect 47762 48628 47768 48680
rect 47820 48668 47826 48680
rect 48593 48671 48651 48677
rect 48593 48668 48605 48671
rect 47820 48640 48605 48668
rect 47820 48628 47826 48640
rect 48593 48637 48605 48640
rect 48639 48637 48651 48671
rect 48593 48631 48651 48637
rect 49099 48671 49157 48677
rect 49099 48637 49111 48671
rect 49145 48668 49157 48671
rect 49234 48668 49240 48680
rect 49145 48640 49240 48668
rect 49145 48637 49157 48640
rect 49099 48631 49157 48637
rect 49234 48628 49240 48640
rect 49292 48628 49298 48680
rect 49326 48628 49332 48680
rect 49384 48668 49390 48680
rect 49384 48640 49429 48668
rect 49384 48628 49390 48640
rect 48038 48600 48044 48612
rect 39908 48572 40080 48600
rect 47999 48572 48044 48600
rect 39908 48560 39914 48572
rect 48038 48560 48044 48572
rect 48096 48560 48102 48612
rect 37550 48492 37556 48544
rect 37608 48532 37614 48544
rect 37737 48535 37795 48541
rect 37737 48532 37749 48535
rect 37608 48504 37749 48532
rect 37608 48492 37614 48504
rect 37737 48501 37749 48504
rect 37783 48532 37795 48535
rect 39482 48532 39488 48544
rect 37783 48504 39488 48532
rect 37783 48501 37795 48504
rect 37737 48495 37795 48501
rect 39482 48492 39488 48504
rect 39540 48492 39546 48544
rect 48133 48535 48191 48541
rect 48133 48501 48145 48535
rect 48179 48532 48191 48535
rect 48406 48532 48412 48544
rect 48179 48504 48412 48532
rect 48179 48501 48191 48504
rect 48133 48495 48191 48501
rect 48406 48492 48412 48504
rect 48464 48492 48470 48544
rect 1104 48442 58880 48464
rect 1104 48390 4214 48442
rect 4266 48390 4278 48442
rect 4330 48390 4342 48442
rect 4394 48390 4406 48442
rect 4458 48390 4470 48442
rect 4522 48390 34934 48442
rect 34986 48390 34998 48442
rect 35050 48390 35062 48442
rect 35114 48390 35126 48442
rect 35178 48390 35190 48442
rect 35242 48390 58880 48442
rect 1104 48368 58880 48390
rect 37458 48328 37464 48340
rect 37419 48300 37464 48328
rect 37458 48288 37464 48300
rect 37516 48288 37522 48340
rect 45002 48288 45008 48340
rect 45060 48328 45066 48340
rect 47762 48328 47768 48340
rect 45060 48300 47768 48328
rect 45060 48288 45066 48300
rect 40129 48195 40187 48201
rect 40129 48161 40141 48195
rect 40175 48192 40187 48195
rect 40218 48192 40224 48204
rect 40175 48164 40224 48192
rect 40175 48161 40187 48164
rect 40129 48155 40187 48161
rect 40218 48152 40224 48164
rect 40276 48152 40282 48204
rect 45664 48192 45692 48300
rect 47762 48288 47768 48300
rect 47820 48288 47826 48340
rect 48130 48288 48136 48340
rect 48188 48328 48194 48340
rect 48225 48331 48283 48337
rect 48225 48328 48237 48331
rect 48188 48300 48237 48328
rect 48188 48288 48194 48300
rect 48225 48297 48237 48300
rect 48271 48297 48283 48331
rect 48225 48291 48283 48297
rect 47581 48263 47639 48269
rect 47581 48229 47593 48263
rect 47627 48260 47639 48263
rect 49326 48260 49332 48272
rect 47627 48232 49332 48260
rect 47627 48229 47639 48232
rect 47581 48223 47639 48229
rect 49326 48220 49332 48232
rect 49384 48220 49390 48272
rect 45741 48195 45799 48201
rect 45741 48192 45753 48195
rect 45664 48164 45753 48192
rect 45741 48161 45753 48164
rect 45787 48161 45799 48195
rect 45741 48155 45799 48161
rect 46014 48152 46020 48204
rect 46072 48192 46078 48204
rect 46204 48195 46262 48201
rect 46204 48192 46216 48195
rect 46072 48164 46216 48192
rect 46072 48152 46078 48164
rect 46204 48161 46216 48164
rect 46250 48161 46262 48195
rect 46204 48155 46262 48161
rect 46382 48152 46388 48204
rect 46440 48192 46446 48204
rect 46477 48195 46535 48201
rect 46477 48192 46489 48195
rect 46440 48164 46489 48192
rect 46440 48152 46446 48164
rect 46477 48161 46489 48164
rect 46523 48192 46535 48195
rect 46842 48192 46848 48204
rect 46523 48164 46848 48192
rect 46523 48161 46535 48164
rect 46477 48155 46535 48161
rect 46842 48152 46848 48164
rect 46900 48152 46906 48204
rect 1946 48084 1952 48136
rect 2004 48124 2010 48136
rect 2041 48127 2099 48133
rect 2041 48124 2053 48127
rect 2004 48096 2053 48124
rect 2004 48084 2010 48096
rect 2041 48093 2053 48096
rect 2087 48093 2099 48127
rect 2041 48087 2099 48093
rect 36722 48084 36728 48136
rect 36780 48124 36786 48136
rect 37185 48127 37243 48133
rect 37185 48124 37197 48127
rect 36780 48096 37197 48124
rect 36780 48084 36786 48096
rect 37185 48093 37197 48096
rect 37231 48124 37243 48127
rect 37826 48124 37832 48136
rect 37231 48096 37832 48124
rect 37231 48093 37243 48096
rect 37185 48087 37243 48093
rect 37826 48084 37832 48096
rect 37884 48084 37890 48136
rect 39298 48084 39304 48136
rect 39356 48124 39362 48136
rect 39853 48127 39911 48133
rect 39853 48124 39865 48127
rect 39356 48096 39865 48124
rect 39356 48084 39362 48096
rect 39853 48093 39865 48096
rect 39899 48124 39911 48127
rect 39942 48124 39948 48136
rect 39899 48096 39948 48124
rect 39899 48093 39911 48096
rect 39853 48087 39911 48093
rect 39942 48084 39948 48096
rect 40000 48084 40006 48136
rect 48406 48124 48412 48136
rect 48367 48096 48412 48124
rect 48406 48084 48412 48096
rect 48464 48084 48470 48136
rect 37461 48059 37519 48065
rect 37461 48025 37473 48059
rect 37507 48056 37519 48059
rect 38562 48056 38568 48068
rect 37507 48028 38568 48056
rect 37507 48025 37519 48028
rect 37461 48019 37519 48025
rect 38562 48016 38568 48028
rect 38620 48016 38626 48068
rect 37277 47991 37335 47997
rect 37277 47957 37289 47991
rect 37323 47988 37335 47991
rect 37366 47988 37372 48000
rect 37323 47960 37372 47988
rect 37323 47957 37335 47960
rect 37277 47951 37335 47957
rect 37366 47948 37372 47960
rect 37424 47948 37430 48000
rect 46198 47948 46204 48000
rect 46256 47997 46262 48000
rect 46256 47988 46265 47997
rect 46256 47960 46301 47988
rect 46256 47951 46265 47960
rect 46256 47948 46262 47951
rect 1104 47898 58880 47920
rect 1104 47846 19574 47898
rect 19626 47846 19638 47898
rect 19690 47846 19702 47898
rect 19754 47846 19766 47898
rect 19818 47846 19830 47898
rect 19882 47846 50294 47898
rect 50346 47846 50358 47898
rect 50410 47846 50422 47898
rect 50474 47846 50486 47898
rect 50538 47846 50550 47898
rect 50602 47846 58880 47898
rect 1104 47824 58880 47846
rect 40310 47744 40316 47796
rect 40368 47784 40374 47796
rect 40503 47787 40561 47793
rect 40503 47784 40515 47787
rect 40368 47756 40515 47784
rect 40368 47744 40374 47756
rect 40503 47753 40515 47756
rect 40549 47784 40561 47787
rect 41046 47784 41052 47796
rect 40549 47756 41052 47784
rect 40549 47753 40561 47756
rect 40503 47747 40561 47753
rect 41046 47744 41052 47756
rect 41104 47744 41110 47796
rect 41598 47744 41604 47796
rect 41656 47784 41662 47796
rect 41877 47787 41935 47793
rect 41877 47784 41889 47787
rect 41656 47756 41889 47784
rect 41656 47744 41662 47756
rect 41877 47753 41889 47756
rect 41923 47753 41935 47787
rect 41877 47747 41935 47753
rect 45649 47787 45707 47793
rect 45649 47753 45661 47787
rect 45695 47784 45707 47787
rect 47670 47784 47676 47796
rect 45695 47756 47676 47784
rect 45695 47753 45707 47756
rect 45649 47747 45707 47753
rect 47670 47744 47676 47756
rect 47728 47744 47734 47796
rect 36633 47719 36691 47725
rect 36633 47685 36645 47719
rect 36679 47716 36691 47719
rect 36679 47688 37412 47716
rect 36679 47685 36691 47688
rect 36633 47679 36691 47685
rect 37384 47660 37412 47688
rect 44726 47676 44732 47728
rect 44784 47716 44790 47728
rect 44784 47688 46704 47716
rect 44784 47676 44790 47688
rect 1946 47648 1952 47660
rect 1907 47620 1952 47648
rect 1946 47608 1952 47620
rect 2004 47608 2010 47660
rect 36357 47651 36415 47657
rect 36357 47617 36369 47651
rect 36403 47648 36415 47651
rect 36446 47648 36452 47660
rect 36403 47620 36452 47648
rect 36403 47617 36415 47620
rect 36357 47611 36415 47617
rect 36446 47608 36452 47620
rect 36504 47608 36510 47660
rect 36722 47648 36728 47660
rect 36683 47620 36728 47648
rect 36722 47608 36728 47620
rect 36780 47608 36786 47660
rect 37366 47608 37372 47660
rect 37424 47648 37430 47660
rect 37737 47651 37795 47657
rect 37737 47648 37749 47651
rect 37424 47620 37749 47648
rect 37424 47608 37430 47620
rect 37737 47617 37749 47620
rect 37783 47617 37795 47651
rect 37737 47611 37795 47617
rect 38562 47608 38568 47660
rect 38620 47648 38626 47660
rect 46382 47648 46388 47660
rect 38620 47620 40356 47648
rect 46343 47620 46388 47648
rect 38620 47608 38626 47620
rect 2133 47583 2191 47589
rect 2133 47549 2145 47583
rect 2179 47580 2191 47583
rect 2406 47580 2412 47592
rect 2179 47552 2412 47580
rect 2179 47549 2191 47552
rect 2133 47543 2191 47549
rect 2406 47540 2412 47552
rect 2464 47540 2470 47592
rect 2774 47580 2780 47592
rect 2735 47552 2780 47580
rect 2774 47540 2780 47552
rect 2832 47540 2838 47592
rect 37461 47583 37519 47589
rect 37461 47549 37473 47583
rect 37507 47580 37519 47583
rect 37550 47580 37556 47592
rect 37507 47552 37556 47580
rect 37507 47549 37519 47552
rect 37461 47543 37519 47549
rect 37550 47540 37556 47552
rect 37608 47580 37614 47592
rect 38470 47580 38476 47592
rect 37608 47552 38476 47580
rect 37608 47540 37614 47552
rect 38470 47540 38476 47552
rect 38528 47540 38534 47592
rect 40037 47583 40095 47589
rect 40037 47549 40049 47583
rect 40083 47580 40095 47583
rect 40218 47580 40224 47592
rect 40083 47552 40224 47580
rect 40083 47549 40095 47552
rect 40037 47543 40095 47549
rect 40218 47540 40224 47552
rect 40276 47540 40282 47592
rect 40328 47580 40356 47620
rect 46382 47608 46388 47620
rect 46440 47608 46446 47660
rect 46676 47657 46704 47688
rect 46661 47651 46719 47657
rect 46661 47617 46673 47651
rect 46707 47648 46719 47651
rect 50798 47648 50804 47660
rect 46707 47620 50804 47648
rect 46707 47617 46719 47620
rect 46661 47611 46719 47617
rect 50798 47608 50804 47620
rect 50856 47608 50862 47660
rect 40500 47583 40558 47589
rect 40500 47580 40512 47583
rect 40328 47552 40512 47580
rect 40500 47549 40512 47552
rect 40546 47549 40558 47583
rect 40500 47543 40558 47549
rect 40773 47583 40831 47589
rect 40773 47549 40785 47583
rect 40819 47580 40831 47583
rect 41874 47580 41880 47592
rect 40819 47552 41880 47580
rect 40819 47549 40831 47552
rect 40773 47543 40831 47549
rect 41874 47540 41880 47552
rect 41932 47540 41938 47592
rect 36354 47444 36360 47456
rect 36315 47416 36360 47444
rect 36354 47404 36360 47416
rect 36412 47404 36418 47456
rect 36449 47447 36507 47453
rect 36449 47413 36461 47447
rect 36495 47444 36507 47447
rect 38194 47444 38200 47456
rect 36495 47416 38200 47444
rect 36495 47413 36507 47416
rect 36449 47407 36507 47413
rect 38194 47404 38200 47416
rect 38252 47404 38258 47456
rect 1104 47354 58880 47376
rect 1104 47302 4214 47354
rect 4266 47302 4278 47354
rect 4330 47302 4342 47354
rect 4394 47302 4406 47354
rect 4458 47302 4470 47354
rect 4522 47302 34934 47354
rect 34986 47302 34998 47354
rect 35050 47302 35062 47354
rect 35114 47302 35126 47354
rect 35178 47302 35190 47354
rect 35242 47302 58880 47354
rect 1104 47280 58880 47302
rect 2406 47240 2412 47252
rect 2367 47212 2412 47240
rect 2406 47200 2412 47212
rect 2464 47200 2470 47252
rect 38194 47240 38200 47252
rect 38155 47212 38200 47240
rect 38194 47200 38200 47212
rect 38252 47200 38258 47252
rect 39298 47240 39304 47252
rect 39259 47212 39304 47240
rect 39298 47200 39304 47212
rect 39356 47200 39362 47252
rect 44726 47240 44732 47252
rect 43456 47212 44732 47240
rect 36354 47132 36360 47184
rect 36412 47132 36418 47184
rect 36372 47104 36400 47132
rect 38933 47107 38991 47113
rect 38933 47104 38945 47107
rect 36372 47076 36492 47104
rect 2501 47039 2559 47045
rect 2501 47005 2513 47039
rect 2547 47036 2559 47039
rect 2590 47036 2596 47048
rect 2547 47008 2596 47036
rect 2547 47005 2559 47008
rect 2501 46999 2559 47005
rect 2590 46996 2596 47008
rect 2648 47036 2654 47048
rect 8846 47036 8852 47048
rect 2648 47008 8852 47036
rect 2648 46996 2654 47008
rect 8846 46996 8852 47008
rect 8904 46996 8910 47048
rect 36262 46996 36268 47048
rect 36320 47036 36326 47048
rect 36357 47039 36415 47045
rect 36357 47036 36369 47039
rect 36320 47008 36369 47036
rect 36320 46996 36326 47008
rect 36357 47005 36369 47008
rect 36403 47005 36415 47039
rect 36464 47036 36492 47076
rect 38396 47076 38945 47104
rect 36613 47039 36671 47045
rect 36613 47036 36625 47039
rect 36464 47008 36625 47036
rect 36357 46999 36415 47005
rect 36613 47005 36625 47008
rect 36659 47005 36671 47039
rect 36613 46999 36671 47005
rect 37642 46996 37648 47048
rect 37700 47036 37706 47048
rect 38396 47045 38424 47076
rect 38933 47073 38945 47076
rect 38979 47073 38991 47107
rect 40126 47104 40132 47116
rect 40087 47076 40132 47104
rect 38933 47067 38991 47073
rect 40126 47064 40132 47076
rect 40184 47064 40190 47116
rect 42794 47064 42800 47116
rect 42852 47104 42858 47116
rect 43456 47113 43484 47212
rect 44726 47200 44732 47212
rect 44784 47200 44790 47252
rect 51813 47243 51871 47249
rect 51813 47209 51825 47243
rect 51859 47240 51871 47243
rect 52730 47240 52736 47252
rect 51859 47212 52736 47240
rect 51859 47209 51871 47212
rect 51813 47203 51871 47209
rect 52730 47200 52736 47212
rect 52788 47200 52794 47252
rect 57977 47175 58035 47181
rect 57977 47172 57989 47175
rect 55186 47144 57989 47172
rect 43441 47107 43499 47113
rect 43441 47104 43453 47107
rect 42852 47076 43453 47104
rect 42852 47064 42858 47076
rect 43441 47073 43453 47076
rect 43487 47073 43499 47107
rect 50798 47104 50804 47116
rect 50759 47076 50804 47104
rect 43441 47067 43499 47073
rect 50798 47064 50804 47076
rect 50856 47064 50862 47116
rect 52270 47104 52276 47116
rect 52231 47076 52276 47104
rect 52270 47064 52276 47076
rect 52328 47064 52334 47116
rect 52638 47113 52644 47116
rect 52596 47107 52644 47113
rect 52596 47073 52608 47107
rect 52642 47073 52644 47107
rect 52596 47067 52644 47073
rect 52638 47064 52644 47067
rect 52696 47064 52702 47116
rect 52779 47107 52837 47113
rect 52779 47073 52791 47107
rect 52825 47104 52837 47107
rect 52914 47104 52920 47116
rect 52825 47076 52920 47104
rect 52825 47073 52837 47076
rect 52779 47067 52837 47073
rect 52914 47064 52920 47076
rect 52972 47064 52978 47116
rect 53009 47107 53067 47113
rect 53009 47073 53021 47107
rect 53055 47104 53067 47107
rect 55186 47104 55214 47144
rect 57977 47141 57989 47144
rect 58023 47141 58035 47175
rect 57977 47135 58035 47141
rect 53055 47076 55214 47104
rect 53055 47073 53067 47076
rect 53009 47067 53067 47073
rect 38381 47039 38439 47045
rect 38381 47036 38393 47039
rect 37700 47008 38393 47036
rect 37700 46996 37706 47008
rect 38381 47005 38393 47008
rect 38427 47005 38439 47039
rect 38381 46999 38439 47005
rect 38470 46996 38476 47048
rect 38528 47036 38534 47048
rect 39114 47036 39120 47048
rect 38528 47008 38573 47036
rect 39075 47008 39120 47036
rect 38528 46996 38534 47008
rect 39114 46996 39120 47008
rect 39172 46996 39178 47048
rect 39666 46996 39672 47048
rect 39724 47036 39730 47048
rect 39853 47039 39911 47045
rect 39853 47036 39865 47039
rect 39724 47008 39865 47036
rect 39724 46996 39730 47008
rect 39853 47005 39865 47008
rect 39899 47005 39911 47039
rect 39853 46999 39911 47005
rect 42981 47039 43039 47045
rect 42981 47005 42993 47039
rect 43027 47036 43039 47039
rect 43070 47036 43076 47048
rect 43027 47008 43076 47036
rect 43027 47005 43039 47008
rect 42981 46999 43039 47005
rect 43070 46996 43076 47008
rect 43128 46996 43134 47048
rect 43622 46996 43628 47048
rect 43680 47036 43686 47048
rect 43717 47039 43775 47045
rect 43717 47036 43729 47039
rect 43680 47008 43729 47036
rect 43680 46996 43686 47008
rect 43717 47005 43729 47008
rect 43763 47036 43775 47039
rect 44358 47036 44364 47048
rect 43763 47008 44364 47036
rect 43763 47005 43775 47008
rect 43717 46999 43775 47005
rect 44358 46996 44364 47008
rect 44416 46996 44422 47048
rect 51074 47036 51080 47048
rect 50987 47008 51080 47036
rect 51074 46996 51080 47008
rect 51132 47036 51138 47048
rect 58158 47036 58164 47048
rect 51132 47008 54156 47036
rect 58119 47008 58164 47036
rect 51132 46996 51138 47008
rect 38197 46971 38255 46977
rect 38197 46968 38209 46971
rect 37752 46940 38209 46968
rect 37752 46909 37780 46940
rect 38197 46937 38209 46940
rect 38243 46968 38255 46971
rect 39132 46968 39160 46996
rect 38243 46940 39160 46968
rect 38243 46937 38255 46940
rect 38197 46931 38255 46937
rect 37737 46903 37795 46909
rect 37737 46869 37749 46903
rect 37783 46869 37795 46903
rect 44450 46900 44456 46912
rect 44411 46872 44456 46900
rect 37737 46863 37795 46869
rect 44450 46860 44456 46872
rect 44508 46860 44514 46912
rect 54128 46909 54156 47008
rect 58158 46996 58164 47008
rect 58216 46996 58222 47048
rect 54113 46903 54171 46909
rect 54113 46869 54125 46903
rect 54159 46869 54171 46903
rect 54113 46863 54171 46869
rect 1104 46810 58880 46832
rect 1104 46758 19574 46810
rect 19626 46758 19638 46810
rect 19690 46758 19702 46810
rect 19754 46758 19766 46810
rect 19818 46758 19830 46810
rect 19882 46758 50294 46810
rect 50346 46758 50358 46810
rect 50410 46758 50422 46810
rect 50474 46758 50486 46810
rect 50538 46758 50550 46810
rect 50602 46758 58880 46810
rect 1104 46736 58880 46758
rect 40310 46656 40316 46708
rect 40368 46696 40374 46708
rect 40503 46699 40561 46705
rect 40503 46696 40515 46699
rect 40368 46668 40515 46696
rect 40368 46656 40374 46668
rect 40503 46665 40515 46668
rect 40549 46696 40561 46699
rect 41874 46696 41880 46708
rect 40549 46668 41736 46696
rect 41835 46668 41880 46696
rect 40549 46665 40561 46668
rect 40503 46659 40561 46665
rect 37369 46631 37427 46637
rect 37369 46597 37381 46631
rect 37415 46628 37427 46631
rect 37642 46628 37648 46640
rect 37415 46600 37648 46628
rect 37415 46597 37427 46600
rect 37369 46591 37427 46597
rect 37642 46588 37648 46600
rect 37700 46588 37706 46640
rect 37277 46563 37335 46569
rect 37277 46529 37289 46563
rect 37323 46529 37335 46563
rect 37277 46523 37335 46529
rect 37553 46563 37611 46569
rect 37553 46529 37565 46563
rect 37599 46560 37611 46563
rect 38654 46560 38660 46572
rect 37599 46532 38660 46560
rect 37599 46529 37611 46532
rect 37553 46523 37611 46529
rect 37292 46424 37320 46523
rect 38654 46520 38660 46532
rect 38712 46520 38718 46572
rect 39114 46520 39120 46572
rect 39172 46560 39178 46572
rect 41708 46560 41736 46668
rect 41874 46656 41880 46668
rect 41932 46656 41938 46708
rect 44358 46656 44364 46708
rect 44416 46696 44422 46708
rect 44453 46699 44511 46705
rect 44453 46696 44465 46699
rect 44416 46668 44465 46696
rect 44416 46656 44422 46668
rect 44453 46665 44465 46668
rect 44499 46665 44511 46699
rect 44453 46659 44511 46665
rect 46198 46656 46204 46708
rect 46256 46696 46262 46708
rect 48038 46696 48044 46708
rect 46256 46668 48044 46696
rect 46256 46656 46262 46668
rect 48038 46656 48044 46668
rect 48096 46696 48102 46708
rect 48954 46699 49012 46705
rect 48954 46696 48966 46699
rect 48096 46668 48966 46696
rect 48096 46656 48102 46668
rect 48954 46665 48966 46668
rect 49000 46696 49012 46699
rect 49418 46696 49424 46708
rect 49000 46668 49424 46696
rect 49000 46665 49012 46668
rect 48954 46659 49012 46665
rect 49418 46656 49424 46668
rect 49476 46656 49482 46708
rect 52733 46699 52791 46705
rect 52733 46665 52745 46699
rect 52779 46665 52791 46699
rect 52733 46659 52791 46665
rect 42936 46563 42994 46569
rect 42936 46560 42948 46563
rect 39172 46532 40172 46560
rect 41708 46532 42948 46560
rect 39172 46520 39178 46532
rect 40037 46495 40095 46501
rect 40037 46461 40049 46495
rect 40083 46461 40095 46495
rect 40144 46492 40172 46532
rect 42936 46529 42948 46532
rect 42982 46560 42994 46563
rect 46198 46560 46204 46572
rect 42982 46532 46204 46560
rect 42982 46529 42994 46532
rect 42936 46523 42994 46529
rect 46198 46520 46204 46532
rect 46256 46520 46262 46572
rect 48685 46563 48743 46569
rect 48685 46529 48697 46563
rect 48731 46560 48743 46563
rect 49602 46560 49608 46572
rect 48731 46532 49608 46560
rect 48731 46529 48743 46532
rect 48685 46523 48743 46529
rect 49602 46520 49608 46532
rect 49660 46520 49666 46572
rect 51169 46563 51227 46569
rect 51169 46529 51181 46563
rect 51215 46560 51227 46563
rect 52748 46560 52776 46659
rect 52917 46631 52975 46637
rect 52917 46597 52929 46631
rect 52963 46628 52975 46631
rect 53006 46628 53012 46640
rect 52963 46600 53012 46628
rect 52963 46597 52975 46600
rect 52917 46591 52975 46597
rect 53006 46588 53012 46600
rect 53064 46588 53070 46640
rect 51215 46532 52776 46560
rect 51215 46529 51227 46532
rect 51169 46523 51227 46529
rect 40500 46513 40558 46519
rect 40500 46492 40512 46513
rect 40144 46479 40512 46492
rect 40546 46479 40558 46513
rect 40144 46473 40558 46479
rect 40773 46495 40831 46501
rect 40144 46464 40540 46473
rect 40037 46455 40095 46461
rect 40773 46461 40785 46495
rect 40819 46492 40831 46495
rect 41782 46492 41788 46504
rect 40819 46464 41788 46492
rect 40819 46461 40831 46464
rect 40773 46455 40831 46461
rect 37366 46424 37372 46436
rect 37292 46396 37372 46424
rect 37366 46384 37372 46396
rect 37424 46384 37430 46436
rect 37458 46316 37464 46368
rect 37516 46356 37522 46368
rect 37553 46359 37611 46365
rect 37553 46356 37565 46359
rect 37516 46328 37565 46356
rect 37516 46316 37522 46328
rect 37553 46325 37565 46328
rect 37599 46325 37611 46359
rect 37553 46319 37611 46325
rect 39850 46316 39856 46368
rect 39908 46356 39914 46368
rect 40052 46356 40080 46455
rect 41782 46452 41788 46464
rect 41840 46452 41846 46504
rect 42334 46452 42340 46504
rect 42392 46492 42398 46504
rect 42613 46495 42671 46501
rect 42613 46492 42625 46495
rect 42392 46464 42625 46492
rect 42392 46452 42398 46464
rect 42613 46461 42625 46464
rect 42659 46461 42671 46495
rect 42613 46455 42671 46461
rect 43070 46452 43076 46504
rect 43128 46492 43134 46504
rect 43349 46495 43407 46501
rect 43128 46464 43173 46492
rect 43128 46452 43134 46464
rect 43349 46461 43361 46495
rect 43395 46492 43407 46495
rect 43395 46464 44220 46492
rect 43395 46461 43407 46464
rect 43349 46455 43407 46461
rect 40218 46356 40224 46368
rect 39908 46328 40224 46356
rect 39908 46316 39914 46328
rect 40218 46316 40224 46328
rect 40276 46356 40282 46368
rect 42352 46356 42380 46452
rect 44192 46436 44220 46464
rect 47026 46452 47032 46504
rect 47084 46492 47090 46504
rect 48915 46495 48973 46501
rect 48915 46492 48927 46495
rect 47084 46464 48927 46492
rect 47084 46452 47090 46464
rect 48915 46461 48927 46464
rect 48961 46461 48973 46495
rect 48915 46455 48973 46461
rect 49421 46495 49479 46501
rect 49421 46461 49433 46495
rect 49467 46461 49479 46495
rect 49421 46455 49479 46461
rect 44174 46384 44180 46436
rect 44232 46424 44238 46436
rect 47581 46427 47639 46433
rect 47581 46424 47593 46427
rect 44232 46396 47593 46424
rect 44232 46384 44238 46396
rect 47581 46393 47593 46396
rect 47627 46393 47639 46427
rect 47581 46387 47639 46393
rect 49436 46424 49464 46455
rect 50798 46424 50804 46436
rect 49436 46396 50804 46424
rect 40276 46328 42380 46356
rect 40276 46316 40282 46328
rect 47762 46316 47768 46368
rect 47820 46356 47826 46368
rect 49436 46356 49464 46396
rect 50798 46384 50804 46396
rect 50856 46384 50862 46436
rect 53282 46424 53288 46436
rect 53243 46396 53288 46424
rect 53282 46384 53288 46396
rect 53340 46384 53346 46436
rect 47820 46328 49464 46356
rect 47820 46316 47826 46328
rect 50614 46316 50620 46368
rect 50672 46356 50678 46368
rect 50985 46359 51043 46365
rect 50985 46356 50997 46359
rect 50672 46328 50997 46356
rect 50672 46316 50678 46328
rect 50985 46325 50997 46328
rect 51031 46325 51043 46359
rect 50985 46319 51043 46325
rect 52730 46316 52736 46368
rect 52788 46356 52794 46368
rect 52917 46359 52975 46365
rect 52917 46356 52929 46359
rect 52788 46328 52929 46356
rect 52788 46316 52794 46328
rect 52917 46325 52929 46328
rect 52963 46325 52975 46359
rect 52917 46319 52975 46325
rect 1104 46266 58880 46288
rect 1104 46214 4214 46266
rect 4266 46214 4278 46266
rect 4330 46214 4342 46266
rect 4394 46214 4406 46266
rect 4458 46214 4470 46266
rect 4522 46214 34934 46266
rect 34986 46214 34998 46266
rect 35050 46214 35062 46266
rect 35114 46214 35126 46266
rect 35178 46214 35190 46266
rect 35242 46214 58880 46266
rect 1104 46192 58880 46214
rect 52089 46087 52147 46093
rect 52089 46053 52101 46087
rect 52135 46084 52147 46087
rect 53282 46084 53288 46096
rect 52135 46056 53288 46084
rect 52135 46053 52147 46056
rect 52089 46047 52147 46053
rect 53282 46044 53288 46056
rect 53340 46044 53346 46096
rect 36262 46016 36268 46028
rect 36223 45988 36268 46016
rect 36262 45976 36268 45988
rect 36320 45976 36326 46028
rect 38105 46019 38163 46025
rect 38105 45985 38117 46019
rect 38151 46016 38163 46019
rect 38654 46016 38660 46028
rect 38151 45988 38660 46016
rect 38151 45985 38163 45988
rect 38105 45979 38163 45985
rect 38654 45976 38660 45988
rect 38712 46016 38718 46028
rect 40126 46016 40132 46028
rect 38712 45988 40132 46016
rect 38712 45976 38718 45988
rect 40126 45976 40132 45988
rect 40184 45976 40190 46028
rect 44453 46019 44511 46025
rect 44453 45985 44465 46019
rect 44499 46016 44511 46019
rect 44726 46016 44732 46028
rect 44499 45988 44732 46016
rect 44499 45985 44511 45988
rect 44453 45979 44511 45985
rect 44726 45976 44732 45988
rect 44784 45976 44790 46028
rect 47762 46016 47768 46028
rect 47723 45988 47768 46016
rect 47762 45976 47768 45988
rect 47820 45976 47826 46028
rect 48038 45976 48044 46028
rect 48096 46025 48102 46028
rect 48096 46019 48146 46025
rect 48096 45985 48100 46019
rect 48134 45985 48146 46019
rect 48096 45979 48146 45985
rect 48096 45976 48102 45979
rect 48222 45976 48228 46028
rect 48280 46016 48286 46028
rect 50982 46016 50988 46028
rect 48280 45988 50988 46016
rect 48280 45976 48286 45988
rect 50982 45976 50988 45988
rect 51040 45976 51046 46028
rect 52914 45976 52920 46028
rect 52972 46016 52978 46028
rect 53009 46019 53067 46025
rect 53009 46016 53021 46019
rect 52972 45988 53021 46016
rect 52972 45976 52978 45988
rect 53009 45985 53021 45988
rect 53055 46016 53067 46019
rect 53190 46016 53196 46028
rect 53055 45988 53196 46016
rect 53055 45985 53067 45988
rect 53009 45979 53067 45985
rect 53190 45976 53196 45988
rect 53248 45976 53254 46028
rect 36354 45908 36360 45960
rect 36412 45948 36418 45960
rect 38381 45951 38439 45957
rect 38381 45948 38393 45951
rect 36412 45920 38393 45948
rect 36412 45908 36418 45920
rect 38381 45917 38393 45920
rect 38427 45917 38439 45951
rect 44174 45948 44180 45960
rect 44135 45920 44180 45948
rect 38381 45911 38439 45917
rect 44174 45908 44180 45920
rect 44232 45908 44238 45960
rect 45649 45951 45707 45957
rect 45649 45917 45661 45951
rect 45695 45917 45707 45951
rect 45649 45911 45707 45917
rect 48501 45951 48559 45957
rect 48501 45917 48513 45951
rect 48547 45948 48559 45951
rect 48547 45920 49280 45948
rect 48547 45917 48559 45920
rect 48501 45911 48559 45917
rect 36532 45883 36590 45889
rect 36532 45849 36544 45883
rect 36578 45880 36590 45883
rect 37274 45880 37280 45892
rect 36578 45852 37280 45880
rect 36578 45849 36590 45852
rect 36532 45843 36590 45849
rect 37274 45840 37280 45852
rect 37332 45840 37338 45892
rect 45664 45880 45692 45911
rect 49252 45892 49280 45920
rect 50890 45908 50896 45960
rect 50948 45948 50954 45960
rect 51077 45951 51135 45957
rect 51077 45948 51089 45951
rect 50948 45920 51089 45948
rect 50948 45908 50954 45920
rect 51077 45917 51089 45920
rect 51123 45917 51135 45951
rect 51077 45911 51135 45917
rect 51353 45951 51411 45957
rect 51353 45917 51365 45951
rect 51399 45917 51411 45951
rect 52730 45948 52736 45960
rect 52691 45920 52736 45948
rect 51353 45911 51411 45917
rect 45922 45889 45928 45892
rect 43456 45852 45692 45880
rect 37642 45812 37648 45824
rect 37603 45784 37648 45812
rect 37642 45772 37648 45784
rect 37700 45772 37706 45824
rect 43070 45772 43076 45824
rect 43128 45812 43134 45824
rect 43456 45821 43484 45852
rect 45916 45843 45928 45889
rect 45980 45880 45986 45892
rect 45980 45852 46016 45880
rect 45922 45840 45928 45843
rect 45980 45840 45986 45852
rect 49234 45840 49240 45892
rect 49292 45880 49298 45892
rect 51368 45880 51396 45911
rect 52730 45908 52736 45920
rect 52788 45908 52794 45960
rect 49292 45852 51396 45880
rect 49292 45840 49298 45852
rect 43441 45815 43499 45821
rect 43441 45812 43453 45815
rect 43128 45784 43453 45812
rect 43128 45772 43134 45784
rect 43441 45781 43453 45784
rect 43487 45781 43499 45815
rect 43441 45775 43499 45781
rect 47029 45815 47087 45821
rect 47029 45781 47041 45815
rect 47075 45812 47087 45815
rect 47118 45812 47124 45824
rect 47075 45784 47124 45812
rect 47075 45781 47087 45784
rect 47029 45775 47087 45781
rect 47118 45772 47124 45784
rect 47176 45812 47182 45824
rect 48038 45812 48044 45824
rect 47176 45784 48044 45812
rect 47176 45772 47182 45784
rect 48038 45772 48044 45784
rect 48096 45772 48102 45824
rect 49605 45815 49663 45821
rect 49605 45781 49617 45815
rect 49651 45812 49663 45815
rect 49878 45812 49884 45824
rect 49651 45784 49884 45812
rect 49651 45781 49663 45784
rect 49605 45775 49663 45781
rect 49878 45772 49884 45784
rect 49936 45772 49942 45824
rect 1104 45722 58880 45744
rect 1104 45670 19574 45722
rect 19626 45670 19638 45722
rect 19690 45670 19702 45722
rect 19754 45670 19766 45722
rect 19818 45670 19830 45722
rect 19882 45670 50294 45722
rect 50346 45670 50358 45722
rect 50410 45670 50422 45722
rect 50474 45670 50486 45722
rect 50538 45670 50550 45722
rect 50602 45670 58880 45722
rect 1104 45648 58880 45670
rect 40310 45568 40316 45620
rect 40368 45608 40374 45620
rect 40411 45611 40469 45617
rect 40411 45608 40423 45611
rect 40368 45580 40423 45608
rect 40368 45568 40374 45580
rect 40411 45577 40423 45580
rect 40457 45577 40469 45611
rect 41782 45608 41788 45620
rect 41743 45580 41788 45608
rect 40411 45571 40469 45577
rect 41782 45568 41788 45580
rect 41840 45568 41846 45620
rect 48961 45611 49019 45617
rect 48961 45577 48973 45611
rect 49007 45608 49019 45611
rect 49234 45608 49240 45620
rect 49007 45580 49240 45608
rect 49007 45577 49019 45580
rect 48961 45571 49019 45577
rect 49234 45568 49240 45580
rect 49292 45568 49298 45620
rect 49418 45568 49424 45620
rect 49476 45608 49482 45620
rect 50334 45611 50392 45617
rect 50334 45608 50346 45611
rect 49476 45580 50346 45608
rect 49476 45568 49482 45580
rect 50334 45577 50346 45580
rect 50380 45577 50392 45611
rect 52730 45608 52736 45620
rect 52691 45580 52736 45608
rect 50334 45571 50392 45577
rect 52730 45568 52736 45580
rect 52788 45568 52794 45620
rect 52917 45611 52975 45617
rect 52917 45577 52929 45611
rect 52963 45608 52975 45611
rect 53282 45608 53288 45620
rect 52963 45580 53288 45608
rect 52963 45577 52975 45580
rect 52917 45571 52975 45577
rect 53282 45568 53288 45580
rect 53340 45568 53346 45620
rect 37274 45540 37280 45552
rect 37235 45512 37280 45540
rect 37274 45500 37280 45512
rect 37332 45500 37338 45552
rect 46845 45543 46903 45549
rect 46845 45509 46857 45543
rect 46891 45540 46903 45543
rect 47026 45540 47032 45552
rect 46891 45512 47032 45540
rect 46891 45509 46903 45512
rect 46845 45503 46903 45509
rect 47026 45500 47032 45512
rect 47084 45500 47090 45552
rect 37458 45472 37464 45484
rect 37419 45444 37464 45472
rect 37458 45432 37464 45444
rect 37516 45432 37522 45484
rect 37642 45432 37648 45484
rect 37700 45472 37706 45484
rect 37737 45475 37795 45481
rect 37737 45472 37749 45475
rect 37700 45444 37749 45472
rect 37700 45432 37706 45444
rect 37737 45441 37749 45444
rect 37783 45472 37795 45475
rect 37783 45444 40356 45472
rect 37783 45441 37795 45444
rect 37737 45435 37795 45441
rect 40328 45422 40356 45444
rect 44174 45432 44180 45484
rect 44232 45472 44238 45484
rect 44361 45475 44419 45481
rect 44361 45472 44373 45475
rect 44232 45444 44373 45472
rect 44232 45432 44238 45444
rect 44361 45441 44373 45444
rect 44407 45441 44419 45475
rect 44361 45435 44419 45441
rect 44450 45432 44456 45484
rect 44508 45472 44514 45484
rect 45097 45475 45155 45481
rect 45097 45472 45109 45475
rect 44508 45444 45109 45472
rect 44508 45432 44514 45444
rect 45097 45441 45109 45444
rect 45143 45441 45155 45475
rect 45554 45472 45560 45484
rect 45515 45444 45560 45472
rect 45097 45435 45155 45441
rect 45554 45432 45560 45444
rect 45612 45432 45618 45484
rect 45833 45475 45891 45481
rect 45833 45441 45845 45475
rect 45879 45472 45891 45475
rect 46477 45475 46535 45481
rect 46477 45472 46489 45475
rect 45879 45444 46489 45472
rect 45879 45441 45891 45444
rect 45833 45435 45891 45441
rect 46477 45441 46489 45444
rect 46523 45441 46535 45475
rect 46477 45435 46535 45441
rect 46937 45475 46995 45481
rect 46937 45441 46949 45475
rect 46983 45472 46995 45475
rect 47394 45472 47400 45484
rect 46983 45444 47400 45472
rect 46983 45441 46995 45444
rect 46937 45435 46995 45441
rect 40408 45425 40466 45431
rect 40408 45422 40420 45425
rect 39850 45364 39856 45416
rect 39908 45404 39914 45416
rect 39945 45407 40003 45413
rect 39945 45404 39957 45407
rect 39908 45376 39957 45404
rect 39908 45364 39914 45376
rect 39945 45373 39957 45376
rect 39991 45373 40003 45407
rect 40328 45394 40420 45422
rect 40408 45391 40420 45394
rect 40454 45391 40466 45425
rect 40408 45385 40466 45391
rect 40681 45407 40739 45413
rect 39945 45367 40003 45373
rect 40681 45373 40693 45407
rect 40727 45404 40739 45407
rect 41690 45404 41696 45416
rect 40727 45376 41696 45404
rect 40727 45373 40739 45376
rect 40681 45367 40739 45373
rect 41690 45364 41696 45376
rect 41748 45364 41754 45416
rect 45462 45404 45468 45416
rect 45423 45376 45468 45404
rect 45462 45364 45468 45376
rect 45520 45364 45526 45416
rect 46492 45404 46520 45435
rect 47394 45432 47400 45444
rect 47452 45432 47458 45484
rect 50065 45475 50123 45481
rect 50065 45441 50077 45475
rect 50111 45472 50123 45475
rect 50111 45444 51074 45472
rect 50111 45441 50123 45444
rect 50065 45435 50123 45441
rect 51046 45416 51074 45444
rect 52822 45432 52828 45484
rect 52880 45472 52886 45484
rect 53285 45475 53343 45481
rect 53285 45472 53297 45475
rect 52880 45444 53297 45472
rect 52880 45432 52886 45444
rect 53285 45441 53297 45444
rect 53331 45441 53343 45475
rect 53285 45435 53343 45441
rect 47118 45404 47124 45416
rect 46492 45376 47124 45404
rect 47118 45364 47124 45376
rect 47176 45364 47182 45416
rect 50295 45407 50353 45413
rect 50295 45373 50307 45407
rect 50341 45404 50353 45407
rect 50614 45404 50620 45416
rect 50341 45376 50620 45404
rect 50341 45373 50353 45376
rect 50295 45367 50353 45373
rect 50614 45364 50620 45376
rect 50672 45364 50678 45416
rect 50798 45404 50804 45416
rect 50759 45376 50804 45404
rect 50798 45364 50804 45376
rect 50856 45364 50862 45416
rect 51046 45376 51080 45416
rect 51074 45364 51080 45376
rect 51132 45364 51138 45416
rect 1946 45228 1952 45280
rect 2004 45268 2010 45280
rect 2041 45271 2099 45277
rect 2041 45268 2053 45271
rect 2004 45240 2053 45268
rect 2004 45228 2010 45240
rect 2041 45237 2053 45240
rect 2087 45237 2099 45271
rect 2041 45231 2099 45237
rect 37366 45228 37372 45280
rect 37424 45268 37430 45280
rect 37645 45271 37703 45277
rect 37645 45268 37657 45271
rect 37424 45240 37657 45268
rect 37424 45228 37430 45240
rect 37645 45237 37657 45240
rect 37691 45237 37703 45271
rect 43898 45268 43904 45280
rect 43859 45240 43904 45268
rect 37645 45231 37703 45237
rect 43898 45228 43904 45240
rect 43956 45228 43962 45280
rect 44269 45271 44327 45277
rect 44269 45237 44281 45271
rect 44315 45268 44327 45271
rect 44450 45268 44456 45280
rect 44315 45240 44456 45268
rect 44315 45237 44327 45240
rect 44269 45231 44327 45237
rect 44450 45228 44456 45240
rect 44508 45228 44514 45280
rect 46658 45277 46664 45280
rect 46615 45271 46664 45277
rect 46615 45237 46627 45271
rect 46661 45237 46664 45271
rect 46615 45231 46664 45237
rect 46658 45228 46664 45231
rect 46716 45228 46722 45280
rect 46750 45228 46756 45280
rect 46808 45268 46814 45280
rect 52917 45271 52975 45277
rect 46808 45240 46853 45268
rect 46808 45228 46814 45240
rect 52917 45237 52929 45271
rect 52963 45268 52975 45271
rect 53006 45268 53012 45280
rect 52963 45240 53012 45268
rect 52963 45237 52975 45240
rect 52917 45231 52975 45237
rect 53006 45228 53012 45240
rect 53064 45228 53070 45280
rect 1104 45178 58880 45200
rect 1104 45126 4214 45178
rect 4266 45126 4278 45178
rect 4330 45126 4342 45178
rect 4394 45126 4406 45178
rect 4458 45126 4470 45178
rect 4522 45126 34934 45178
rect 34986 45126 34998 45178
rect 35050 45126 35062 45178
rect 35114 45126 35126 45178
rect 35178 45126 35190 45178
rect 35242 45126 58880 45178
rect 1104 45104 58880 45126
rect 41690 45064 41696 45076
rect 41651 45036 41696 45064
rect 41690 45024 41696 45036
rect 41748 45024 41754 45076
rect 45833 45067 45891 45073
rect 45833 45033 45845 45067
rect 45879 45064 45891 45067
rect 45922 45064 45928 45076
rect 45879 45036 45928 45064
rect 45879 45033 45891 45036
rect 45833 45027 45891 45033
rect 45922 45024 45928 45036
rect 45980 45024 45986 45076
rect 46658 45024 46664 45076
rect 46716 45064 46722 45076
rect 46937 45067 46995 45073
rect 46937 45064 46949 45067
rect 46716 45036 46949 45064
rect 46716 45024 46722 45036
rect 46937 45033 46949 45036
rect 46983 45033 46995 45067
rect 47394 45064 47400 45076
rect 47355 45036 47400 45064
rect 46937 45027 46995 45033
rect 47394 45024 47400 45036
rect 47452 45024 47458 45076
rect 47581 45067 47639 45073
rect 47581 45033 47593 45067
rect 47627 45033 47639 45067
rect 50890 45064 50896 45076
rect 47581 45027 47639 45033
rect 50448 45036 50896 45064
rect 36909 44999 36967 45005
rect 36909 44965 36921 44999
rect 36955 44996 36967 44999
rect 37737 44999 37795 45005
rect 37737 44996 37749 44999
rect 36955 44968 37749 44996
rect 36955 44965 36967 44968
rect 36909 44959 36967 44965
rect 37737 44965 37749 44968
rect 37783 44965 37795 44999
rect 37737 44959 37795 44965
rect 36446 44888 36452 44940
rect 36504 44928 36510 44940
rect 36725 44931 36783 44937
rect 36725 44928 36737 44931
rect 36504 44900 36737 44928
rect 36504 44888 36510 44900
rect 36725 44897 36737 44900
rect 36771 44897 36783 44931
rect 36725 44891 36783 44897
rect 39482 44888 39488 44940
rect 39540 44928 39546 44940
rect 40316 44931 40374 44937
rect 40316 44928 40328 44931
rect 39540 44900 40328 44928
rect 39540 44888 39546 44900
rect 40316 44897 40328 44900
rect 40362 44897 40374 44931
rect 40316 44891 40374 44897
rect 45462 44888 45468 44940
rect 45520 44928 45526 44940
rect 46934 44928 46940 44940
rect 45520 44900 45692 44928
rect 45520 44888 45526 44900
rect 2498 44860 2504 44872
rect 2459 44832 2504 44860
rect 2498 44820 2504 44832
rect 2556 44820 2562 44872
rect 37001 44863 37059 44869
rect 37001 44829 37013 44863
rect 37047 44860 37059 44863
rect 37366 44860 37372 44872
rect 37047 44832 37372 44860
rect 37047 44829 37059 44832
rect 37001 44823 37059 44829
rect 37366 44820 37372 44832
rect 37424 44820 37430 44872
rect 37458 44820 37464 44872
rect 37516 44860 37522 44872
rect 37737 44863 37795 44869
rect 37516 44832 37561 44860
rect 37516 44820 37522 44832
rect 37737 44829 37749 44863
rect 37783 44860 37795 44863
rect 39500 44860 39528 44888
rect 39850 44860 39856 44872
rect 37783 44832 39528 44860
rect 39811 44832 39856 44860
rect 37783 44829 37795 44832
rect 37737 44823 37795 44829
rect 39850 44820 39856 44832
rect 39908 44820 39914 44872
rect 40589 44863 40647 44869
rect 40589 44829 40601 44863
rect 40635 44860 40647 44863
rect 41690 44860 41696 44872
rect 40635 44832 41696 44860
rect 40635 44829 40647 44832
rect 40589 44823 40647 44829
rect 41690 44820 41696 44832
rect 41748 44820 41754 44872
rect 43070 44860 43076 44872
rect 43031 44832 43076 44860
rect 43070 44820 43076 44832
rect 43128 44820 43134 44872
rect 45373 44863 45431 44869
rect 45373 44829 45385 44863
rect 45419 44860 45431 44863
rect 45554 44860 45560 44872
rect 45419 44832 45560 44860
rect 45419 44829 45431 44832
rect 45373 44823 45431 44829
rect 45554 44820 45560 44832
rect 45612 44820 45618 44872
rect 45664 44869 45692 44900
rect 46492 44900 46940 44928
rect 45649 44863 45707 44869
rect 45649 44829 45661 44863
rect 45695 44829 45707 44863
rect 46290 44860 46296 44872
rect 46251 44832 46296 44860
rect 45649 44823 45707 44829
rect 46290 44820 46296 44832
rect 46348 44820 46354 44872
rect 46492 44869 46520 44900
rect 46934 44888 46940 44900
rect 46992 44928 46998 44940
rect 47596 44928 47624 45027
rect 46992 44900 47624 44928
rect 46992 44888 46998 44900
rect 50154 44888 50160 44940
rect 50212 44928 50218 44940
rect 50448 44937 50476 45036
rect 50890 45024 50896 45036
rect 50948 45064 50954 45076
rect 50948 45036 51948 45064
rect 50948 45024 50954 45036
rect 51920 44937 51948 45036
rect 50433 44931 50491 44937
rect 50433 44928 50445 44931
rect 50212 44900 50445 44928
rect 50212 44888 50218 44900
rect 50433 44897 50445 44900
rect 50479 44897 50491 44931
rect 50433 44891 50491 44897
rect 51905 44931 51963 44937
rect 51905 44897 51917 44931
rect 51951 44897 51963 44931
rect 51905 44891 51963 44897
rect 46477 44863 46535 44869
rect 46477 44829 46489 44863
rect 46523 44829 46535 44863
rect 46477 44823 46535 44829
rect 46566 44820 46572 44872
rect 46624 44860 46630 44872
rect 46707 44863 46765 44869
rect 46624 44832 46669 44860
rect 46624 44820 46630 44832
rect 46707 44829 46719 44863
rect 46753 44860 46765 44863
rect 46842 44860 46848 44872
rect 46753 44832 46848 44860
rect 46753 44829 46765 44832
rect 46707 44823 46765 44829
rect 46842 44820 46848 44832
rect 46900 44860 46906 44872
rect 47581 44863 47639 44869
rect 47581 44860 47593 44863
rect 46900 44832 47593 44860
rect 46900 44820 46906 44832
rect 47581 44829 47593 44832
rect 47627 44829 47639 44863
rect 47581 44823 47639 44829
rect 47670 44820 47676 44872
rect 47728 44860 47734 44872
rect 48038 44860 48044 44872
rect 47728 44832 47773 44860
rect 47999 44832 48044 44860
rect 47728 44820 47734 44832
rect 48038 44820 48044 44832
rect 48096 44820 48102 44872
rect 49878 44820 49884 44872
rect 49936 44860 49942 44872
rect 50709 44863 50767 44869
rect 50709 44860 50721 44863
rect 49936 44832 50721 44860
rect 49936 44820 49942 44832
rect 50709 44829 50721 44832
rect 50755 44829 50767 44863
rect 50709 44823 50767 44829
rect 52181 44863 52239 44869
rect 52181 44829 52193 44863
rect 52227 44829 52239 44863
rect 52181 44823 52239 44829
rect 43340 44795 43398 44801
rect 43340 44761 43352 44795
rect 43386 44792 43398 44795
rect 43714 44792 43720 44804
rect 43386 44764 43720 44792
rect 43386 44761 43398 44764
rect 43340 44755 43398 44761
rect 43714 44752 43720 44764
rect 43772 44752 43778 44804
rect 45465 44795 45523 44801
rect 45465 44761 45477 44795
rect 45511 44792 45523 44795
rect 47118 44792 47124 44804
rect 45511 44764 47124 44792
rect 45511 44761 45523 44764
rect 45465 44755 45523 44761
rect 47118 44752 47124 44764
rect 47176 44752 47182 44804
rect 52196 44792 52224 44823
rect 52362 44792 52368 44804
rect 52196 44764 52368 44792
rect 52362 44752 52368 44764
rect 52420 44752 52426 44804
rect 2130 44684 2136 44736
rect 2188 44724 2194 44736
rect 2409 44727 2467 44733
rect 2409 44724 2421 44727
rect 2188 44696 2421 44724
rect 2188 44684 2194 44696
rect 2409 44693 2421 44696
rect 2455 44693 2467 44727
rect 36998 44724 37004 44736
rect 36959 44696 37004 44724
rect 2409 44687 2467 44693
rect 36998 44684 37004 44696
rect 37056 44684 37062 44736
rect 37553 44727 37611 44733
rect 37553 44693 37565 44727
rect 37599 44724 37611 44727
rect 38654 44724 38660 44736
rect 37599 44696 38660 44724
rect 37599 44693 37611 44696
rect 37553 44687 37611 44693
rect 38654 44684 38660 44696
rect 38712 44684 38718 44736
rect 40310 44684 40316 44736
rect 40368 44733 40374 44736
rect 40368 44724 40377 44733
rect 44450 44724 44456 44736
rect 40368 44696 40413 44724
rect 44411 44696 44456 44724
rect 40368 44687 40377 44696
rect 40368 44684 40374 44687
rect 44450 44684 44456 44696
rect 44508 44684 44514 44736
rect 51442 44724 51448 44736
rect 51403 44696 51448 44724
rect 51442 44684 51448 44696
rect 51500 44684 51506 44736
rect 52730 44684 52736 44736
rect 52788 44724 52794 44736
rect 52917 44727 52975 44733
rect 52917 44724 52929 44727
rect 52788 44696 52929 44724
rect 52788 44684 52794 44696
rect 52917 44693 52929 44696
rect 52963 44693 52975 44727
rect 52917 44687 52975 44693
rect 1104 44634 58880 44656
rect 1104 44582 19574 44634
rect 19626 44582 19638 44634
rect 19690 44582 19702 44634
rect 19754 44582 19766 44634
rect 19818 44582 19830 44634
rect 19882 44582 50294 44634
rect 50346 44582 50358 44634
rect 50410 44582 50422 44634
rect 50474 44582 50486 44634
rect 50538 44582 50550 44634
rect 50602 44582 58880 44634
rect 1104 44560 58880 44582
rect 38657 44523 38715 44529
rect 38657 44489 38669 44523
rect 38703 44520 38715 44523
rect 39482 44520 39488 44532
rect 39540 44529 39546 44532
rect 39540 44523 39559 44529
rect 38703 44492 39488 44520
rect 38703 44489 38715 44492
rect 38657 44483 38715 44489
rect 39482 44480 39488 44492
rect 39547 44489 39559 44523
rect 39666 44520 39672 44532
rect 39627 44492 39672 44520
rect 39540 44483 39559 44489
rect 39540 44480 39546 44483
rect 39666 44480 39672 44492
rect 39724 44480 39730 44532
rect 40126 44520 40132 44532
rect 40087 44492 40132 44520
rect 40126 44480 40132 44492
rect 40184 44480 40190 44532
rect 43714 44520 43720 44532
rect 43675 44492 43720 44520
rect 43714 44480 43720 44492
rect 43772 44480 43778 44532
rect 49418 44480 49424 44532
rect 49476 44520 49482 44532
rect 49611 44523 49669 44529
rect 49611 44520 49623 44523
rect 49476 44492 49623 44520
rect 49476 44480 49482 44492
rect 49611 44489 49623 44492
rect 49657 44489 49669 44523
rect 53006 44520 53012 44532
rect 52967 44492 53012 44520
rect 49611 44483 49669 44489
rect 53006 44480 53012 44492
rect 53064 44480 53070 44532
rect 2130 44452 2136 44464
rect 2091 44424 2136 44452
rect 2130 44412 2136 44424
rect 2188 44412 2194 44464
rect 36998 44412 37004 44464
rect 37056 44452 37062 44464
rect 37522 44455 37580 44461
rect 37522 44452 37534 44455
rect 37056 44424 37534 44452
rect 37056 44412 37062 44424
rect 37522 44421 37534 44424
rect 37568 44421 37580 44455
rect 37522 44415 37580 44421
rect 39301 44455 39359 44461
rect 39301 44421 39313 44455
rect 39347 44421 39359 44455
rect 46934 44452 46940 44464
rect 39301 44415 39359 44421
rect 46216 44424 46940 44452
rect 1946 44384 1952 44396
rect 1907 44356 1952 44384
rect 1946 44344 1952 44356
rect 2004 44344 2010 44396
rect 36262 44344 36268 44396
rect 36320 44384 36326 44396
rect 37274 44384 37280 44396
rect 36320 44356 37280 44384
rect 36320 44344 36326 44356
rect 37274 44344 37280 44356
rect 37332 44344 37338 44396
rect 38654 44344 38660 44396
rect 38712 44384 38718 44396
rect 39316 44384 39344 44415
rect 38712 44356 39344 44384
rect 40865 44387 40923 44393
rect 38712 44344 38718 44356
rect 40865 44353 40877 44387
rect 40911 44384 40923 44387
rect 41690 44384 41696 44396
rect 40911 44356 41696 44384
rect 40911 44353 40923 44356
rect 40865 44347 40923 44353
rect 41690 44344 41696 44356
rect 41748 44344 41754 44396
rect 43898 44384 43904 44396
rect 43859 44356 43904 44384
rect 43898 44344 43904 44356
rect 43956 44344 43962 44396
rect 44450 44344 44456 44396
rect 44508 44384 44514 44396
rect 44637 44387 44695 44393
rect 44637 44384 44649 44387
rect 44508 44356 44649 44384
rect 44508 44344 44514 44356
rect 44637 44353 44649 44356
rect 44683 44384 44695 44387
rect 45370 44384 45376 44396
rect 44683 44356 45376 44384
rect 44683 44353 44695 44356
rect 44637 44347 44695 44353
rect 45370 44344 45376 44356
rect 45428 44344 45434 44396
rect 46216 44393 46244 44424
rect 46934 44412 46940 44424
rect 46992 44412 46998 44464
rect 52730 44452 52736 44464
rect 52691 44424 52736 44452
rect 52730 44412 52736 44424
rect 52788 44412 52794 44464
rect 46201 44387 46259 44393
rect 46201 44353 46213 44387
rect 46247 44353 46259 44387
rect 46201 44347 46259 44353
rect 46290 44344 46296 44396
rect 46348 44384 46354 44396
rect 46477 44387 46535 44393
rect 46348 44356 46441 44384
rect 46348 44344 46354 44356
rect 46477 44353 46489 44387
rect 46523 44384 46535 44387
rect 46842 44384 46848 44396
rect 46523 44356 46848 44384
rect 46523 44353 46535 44356
rect 46477 44347 46535 44353
rect 2774 44316 2780 44328
rect 2735 44288 2780 44316
rect 2774 44276 2780 44288
rect 2832 44276 2838 44328
rect 41141 44319 41199 44325
rect 41141 44285 41153 44319
rect 41187 44316 41199 44319
rect 41506 44316 41512 44328
rect 41187 44288 41512 44316
rect 41187 44285 41199 44288
rect 41141 44279 41199 44285
rect 41506 44276 41512 44288
rect 41564 44316 41570 44328
rect 42702 44316 42708 44328
rect 41564 44288 42708 44316
rect 41564 44276 41570 44288
rect 42702 44276 42708 44288
rect 42760 44276 42766 44328
rect 44174 44276 44180 44328
rect 44232 44316 44238 44328
rect 44913 44319 44971 44325
rect 44913 44316 44925 44319
rect 44232 44288 44925 44316
rect 44232 44276 44238 44288
rect 44913 44285 44925 44288
rect 44959 44316 44971 44319
rect 46308 44316 46336 44344
rect 46492 44316 46520 44347
rect 46842 44344 46848 44356
rect 46900 44344 46906 44396
rect 49878 44384 49884 44396
rect 49839 44356 49884 44384
rect 49878 44344 49884 44356
rect 49936 44344 49942 44396
rect 53006 44384 53012 44396
rect 52967 44356 53012 44384
rect 53006 44344 53012 44356
rect 53064 44344 53070 44396
rect 49694 44325 49700 44328
rect 44959 44288 46336 44316
rect 46400 44288 46520 44316
rect 49145 44319 49203 44325
rect 44959 44285 44971 44288
rect 44913 44279 44971 44285
rect 45278 44208 45284 44260
rect 45336 44248 45342 44260
rect 46400 44248 46428 44288
rect 49145 44285 49157 44319
rect 49191 44285 49203 44319
rect 49651 44319 49700 44325
rect 49651 44316 49663 44319
rect 49607 44288 49663 44316
rect 49145 44279 49203 44285
rect 49651 44285 49663 44288
rect 49697 44285 49700 44319
rect 49651 44279 49700 44285
rect 45336 44220 46428 44248
rect 46477 44251 46535 44257
rect 45336 44208 45342 44220
rect 46477 44217 46489 44251
rect 46523 44248 46535 44251
rect 46750 44248 46756 44260
rect 46523 44220 46756 44248
rect 46523 44217 46535 44220
rect 46477 44211 46535 44217
rect 46750 44208 46756 44220
rect 46808 44208 46814 44260
rect 39482 44180 39488 44192
rect 39443 44152 39488 44180
rect 39482 44140 39488 44152
rect 39540 44140 39546 44192
rect 49160 44180 49188 44279
rect 49694 44276 49700 44279
rect 49752 44316 49758 44328
rect 50614 44316 50620 44328
rect 49752 44288 50620 44316
rect 49752 44276 49758 44288
rect 50614 44276 50620 44288
rect 50672 44276 50678 44328
rect 51442 44276 51448 44328
rect 51500 44316 51506 44328
rect 52917 44319 52975 44325
rect 52917 44316 52929 44319
rect 51500 44288 52929 44316
rect 51500 44276 51506 44288
rect 52917 44285 52929 44288
rect 52963 44285 52975 44319
rect 52917 44279 52975 44285
rect 50062 44180 50068 44192
rect 49160 44152 50068 44180
rect 50062 44140 50068 44152
rect 50120 44180 50126 44192
rect 50798 44180 50804 44192
rect 50120 44152 50804 44180
rect 50120 44140 50126 44152
rect 50798 44140 50804 44152
rect 50856 44140 50862 44192
rect 50985 44183 51043 44189
rect 50985 44149 50997 44183
rect 51031 44180 51043 44183
rect 52362 44180 52368 44192
rect 51031 44152 52368 44180
rect 51031 44149 51043 44152
rect 50985 44143 51043 44149
rect 52362 44140 52368 44152
rect 52420 44140 52426 44192
rect 1104 44090 58880 44112
rect 1104 44038 4214 44090
rect 4266 44038 4278 44090
rect 4330 44038 4342 44090
rect 4394 44038 4406 44090
rect 4458 44038 4470 44090
rect 4522 44038 34934 44090
rect 34986 44038 34998 44090
rect 35050 44038 35062 44090
rect 35114 44038 35126 44090
rect 35178 44038 35190 44090
rect 35242 44038 58880 44090
rect 1104 44016 58880 44038
rect 37274 43936 37280 43988
rect 37332 43976 37338 43988
rect 40497 43979 40555 43985
rect 40497 43976 40509 43979
rect 37332 43948 40509 43976
rect 37332 43936 37338 43948
rect 40497 43945 40509 43948
rect 40543 43945 40555 43979
rect 40497 43939 40555 43945
rect 46566 43936 46572 43988
rect 46624 43976 46630 43988
rect 46661 43979 46719 43985
rect 46661 43976 46673 43979
rect 46624 43948 46673 43976
rect 46624 43936 46630 43948
rect 46661 43945 46673 43948
rect 46707 43945 46719 43979
rect 46661 43939 46719 43945
rect 36446 43868 36452 43920
rect 36504 43908 36510 43920
rect 37918 43908 37924 43920
rect 36504 43880 37924 43908
rect 36504 43868 36510 43880
rect 37918 43868 37924 43880
rect 37976 43868 37982 43920
rect 38013 43911 38071 43917
rect 38013 43877 38025 43911
rect 38059 43877 38071 43911
rect 38013 43871 38071 43877
rect 38028 43840 38056 43871
rect 37292 43812 38056 43840
rect 37292 43781 37320 43812
rect 41506 43800 41512 43852
rect 41564 43840 41570 43852
rect 41564 43812 41609 43840
rect 41564 43800 41570 43812
rect 37277 43775 37335 43781
rect 37277 43741 37289 43775
rect 37323 43741 37335 43775
rect 37458 43772 37464 43784
rect 37419 43744 37464 43772
rect 37277 43735 37335 43741
rect 37458 43732 37464 43744
rect 37516 43732 37522 43784
rect 37553 43775 37611 43781
rect 37553 43741 37565 43775
rect 37599 43741 37611 43775
rect 37553 43735 37611 43741
rect 36906 43596 36912 43648
rect 36964 43636 36970 43648
rect 37093 43639 37151 43645
rect 37093 43636 37105 43639
rect 36964 43608 37105 43636
rect 36964 43596 36970 43608
rect 37093 43605 37105 43608
rect 37139 43605 37151 43639
rect 37568 43636 37596 43735
rect 37642 43732 37648 43784
rect 37700 43772 37706 43784
rect 38286 43772 38292 43784
rect 37700 43744 38292 43772
rect 37700 43732 37706 43744
rect 38286 43732 38292 43744
rect 38344 43772 38350 43784
rect 39482 43772 39488 43784
rect 38344 43744 39488 43772
rect 38344 43732 38350 43744
rect 39482 43732 39488 43744
rect 39540 43732 39546 43784
rect 40494 43732 40500 43784
rect 40552 43772 40558 43784
rect 41233 43775 41291 43781
rect 41233 43772 41245 43775
rect 40552 43744 41245 43772
rect 40552 43732 40558 43744
rect 41233 43741 41245 43744
rect 41279 43741 41291 43775
rect 41233 43735 41291 43741
rect 44085 43775 44143 43781
rect 44085 43741 44097 43775
rect 44131 43772 44143 43775
rect 44174 43772 44180 43784
rect 44131 43744 44180 43772
rect 44131 43741 44143 43744
rect 44085 43735 44143 43741
rect 44174 43732 44180 43744
rect 44232 43732 44238 43784
rect 44269 43775 44327 43781
rect 44269 43741 44281 43775
rect 44315 43772 44327 43775
rect 45278 43772 45284 43784
rect 44315 43744 45284 43772
rect 44315 43741 44327 43744
rect 44269 43735 44327 43741
rect 45278 43732 45284 43744
rect 45336 43732 45342 43784
rect 46753 43775 46811 43781
rect 46753 43741 46765 43775
rect 46799 43772 46811 43775
rect 47026 43772 47032 43784
rect 46799 43744 47032 43772
rect 46799 43741 46811 43744
rect 46753 43735 46811 43741
rect 47026 43732 47032 43744
rect 47084 43772 47090 43784
rect 47670 43772 47676 43784
rect 47084 43744 47676 43772
rect 47084 43732 47090 43744
rect 47670 43732 47676 43744
rect 47728 43732 47734 43784
rect 37918 43664 37924 43716
rect 37976 43704 37982 43716
rect 38013 43707 38071 43713
rect 38013 43704 38025 43707
rect 37976 43676 38025 43704
rect 37976 43664 37982 43676
rect 38013 43673 38025 43676
rect 38059 43673 38071 43707
rect 38013 43667 38071 43673
rect 38197 43639 38255 43645
rect 38197 43636 38209 43639
rect 37568 43608 38209 43636
rect 37093 43599 37151 43605
rect 38197 43605 38209 43608
rect 38243 43636 38255 43639
rect 38654 43636 38660 43648
rect 38243 43608 38660 43636
rect 38243 43605 38255 43608
rect 38197 43599 38255 43605
rect 38654 43596 38660 43608
rect 38712 43596 38718 43648
rect 44266 43636 44272 43648
rect 44227 43608 44272 43636
rect 44266 43596 44272 43608
rect 44324 43596 44330 43648
rect 1104 43546 58880 43568
rect 1104 43494 19574 43546
rect 19626 43494 19638 43546
rect 19690 43494 19702 43546
rect 19754 43494 19766 43546
rect 19818 43494 19830 43546
rect 19882 43494 50294 43546
rect 50346 43494 50358 43546
rect 50410 43494 50422 43546
rect 50474 43494 50486 43546
rect 50538 43494 50550 43546
rect 50602 43494 58880 43546
rect 1104 43472 58880 43494
rect 40310 43432 40316 43444
rect 40368 43441 40374 43444
rect 40229 43404 40316 43432
rect 40310 43392 40316 43404
rect 40368 43432 40377 43441
rect 41230 43432 41236 43444
rect 40368 43404 41236 43432
rect 40368 43395 40377 43404
rect 40368 43392 40374 43395
rect 41230 43392 41236 43404
rect 41288 43392 41294 43444
rect 41690 43432 41696 43444
rect 41651 43404 41696 43432
rect 41690 43392 41696 43404
rect 41748 43392 41754 43444
rect 45554 43392 45560 43444
rect 45612 43432 45618 43444
rect 45922 43432 45928 43444
rect 45612 43404 45928 43432
rect 45612 43392 45618 43404
rect 45922 43392 45928 43404
rect 45980 43432 45986 43444
rect 46109 43435 46167 43441
rect 46109 43432 46121 43435
rect 45980 43404 46121 43432
rect 45980 43392 45986 43404
rect 46109 43401 46121 43404
rect 46155 43401 46167 43435
rect 46109 43395 46167 43401
rect 49418 43392 49424 43444
rect 49476 43432 49482 43444
rect 49598 43435 49656 43441
rect 49598 43432 49610 43435
rect 49476 43404 49610 43432
rect 49476 43392 49482 43404
rect 49598 43401 49610 43404
rect 49644 43401 49656 43435
rect 49598 43395 49656 43401
rect 53006 43392 53012 43444
rect 53064 43432 53070 43444
rect 53193 43435 53251 43441
rect 53193 43432 53205 43435
rect 53064 43404 53205 43432
rect 53064 43392 53070 43404
rect 53193 43401 53205 43404
rect 53239 43401 53251 43435
rect 53193 43395 53251 43401
rect 36633 43367 36691 43373
rect 36633 43333 36645 43367
rect 36679 43364 36691 43367
rect 37522 43367 37580 43373
rect 37522 43364 37534 43367
rect 36679 43336 37534 43364
rect 36679 43333 36691 43336
rect 36633 43327 36691 43333
rect 37522 43333 37534 43336
rect 37568 43333 37580 43367
rect 37522 43327 37580 43333
rect 43901 43367 43959 43373
rect 43901 43333 43913 43367
rect 43947 43364 43959 43367
rect 44174 43364 44180 43376
rect 43947 43336 44180 43364
rect 43947 43333 43959 43336
rect 43901 43327 43959 43333
rect 44174 43324 44180 43336
rect 44232 43324 44238 43376
rect 46569 43367 46627 43373
rect 46569 43333 46581 43367
rect 46615 43364 46627 43367
rect 47026 43364 47032 43376
rect 46615 43336 47032 43364
rect 46615 43333 46627 43336
rect 46569 43327 46627 43333
rect 47026 43324 47032 43336
rect 47084 43324 47090 43376
rect 36446 43256 36452 43308
rect 36504 43296 36510 43308
rect 36541 43299 36599 43305
rect 36541 43296 36553 43299
rect 36504 43268 36553 43296
rect 36504 43256 36510 43268
rect 36541 43265 36553 43268
rect 36587 43265 36599 43299
rect 36541 43259 36599 43265
rect 36725 43299 36783 43305
rect 36725 43265 36737 43299
rect 36771 43296 36783 43299
rect 38654 43296 38660 43308
rect 36771 43268 38660 43296
rect 36771 43265 36783 43268
rect 36725 43259 36783 43265
rect 38654 43256 38660 43268
rect 38712 43256 38718 43308
rect 39482 43256 39488 43308
rect 39540 43296 39546 43308
rect 44085 43299 44143 43305
rect 39540 43268 39988 43296
rect 39540 43256 39546 43268
rect 37274 43228 37280 43240
rect 37235 43200 37280 43228
rect 37274 43188 37280 43200
rect 37332 43188 37338 43240
rect 39850 43228 39856 43240
rect 39763 43200 39856 43228
rect 39850 43188 39856 43200
rect 39908 43188 39914 43240
rect 39960 43228 39988 43268
rect 44085 43265 44097 43299
rect 44131 43296 44143 43299
rect 45278 43296 45284 43308
rect 44131 43268 45284 43296
rect 44131 43265 44143 43268
rect 44085 43259 44143 43265
rect 45278 43256 45284 43268
rect 45336 43256 45342 43308
rect 46293 43299 46351 43305
rect 46293 43296 46305 43299
rect 45572 43268 46305 43296
rect 40316 43249 40374 43255
rect 40316 43228 40328 43249
rect 39960 43215 40328 43228
rect 40362 43215 40374 43249
rect 45572 43240 45600 43268
rect 46293 43265 46305 43268
rect 46339 43265 46351 43299
rect 46293 43259 46351 43265
rect 52454 43256 52460 43308
rect 52512 43296 52518 43308
rect 52733 43299 52791 43305
rect 52733 43296 52745 43299
rect 52512 43268 52745 43296
rect 52512 43256 52518 43268
rect 52733 43265 52745 43268
rect 52779 43265 52791 43299
rect 52733 43259 52791 43265
rect 52822 43256 52828 43308
rect 52880 43296 52886 43308
rect 53009 43299 53067 43305
rect 53009 43296 53021 43299
rect 52880 43268 53021 43296
rect 52880 43256 52886 43268
rect 53009 43265 53021 43268
rect 53055 43265 53067 43299
rect 53009 43259 53067 43265
rect 49602 43249 49660 43255
rect 39960 43209 40374 43215
rect 39960 43200 40356 43209
rect 40494 43188 40500 43240
rect 40552 43228 40558 43240
rect 40589 43231 40647 43237
rect 40589 43228 40601 43231
rect 40552 43200 40601 43228
rect 40552 43188 40558 43200
rect 40589 43197 40601 43200
rect 40635 43197 40647 43231
rect 45554 43228 45560 43240
rect 45515 43200 45560 43228
rect 40589 43191 40647 43197
rect 45554 43188 45560 43200
rect 45612 43188 45618 43240
rect 46477 43231 46535 43237
rect 46477 43197 46489 43231
rect 46523 43228 46535 43231
rect 46934 43228 46940 43240
rect 46523 43200 46940 43228
rect 46523 43197 46535 43200
rect 46477 43191 46535 43197
rect 46934 43188 46940 43200
rect 46992 43188 46998 43240
rect 49326 43228 49332 43240
rect 49287 43200 49332 43228
rect 49326 43188 49332 43200
rect 49384 43188 49390 43240
rect 49602 43215 49614 43249
rect 49648 43228 49660 43249
rect 49694 43228 49700 43240
rect 49648 43215 49700 43228
rect 49602 43209 49700 43215
rect 49620 43200 49700 43209
rect 49694 43188 49700 43200
rect 49752 43188 49758 43240
rect 50062 43228 50068 43240
rect 50023 43200 50068 43228
rect 50062 43188 50068 43200
rect 50120 43188 50126 43240
rect 52914 43228 52920 43240
rect 52875 43200 52920 43228
rect 52914 43188 52920 43200
rect 52972 43188 52978 43240
rect 2593 43095 2651 43101
rect 2593 43061 2605 43095
rect 2639 43092 2651 43095
rect 4062 43092 4068 43104
rect 2639 43064 4068 43092
rect 2639 43061 2651 43064
rect 2593 43055 2651 43061
rect 4062 43052 4068 43064
rect 4120 43052 4126 43104
rect 38654 43092 38660 43104
rect 38615 43064 38660 43092
rect 38654 43052 38660 43064
rect 38712 43052 38718 43104
rect 39868 43092 39896 43188
rect 53006 43160 53012 43172
rect 51046 43132 53012 43160
rect 41506 43092 41512 43104
rect 39868 43064 41512 43092
rect 41506 43052 41512 43064
rect 41564 43052 41570 43104
rect 44174 43052 44180 43104
rect 44232 43092 44238 43104
rect 44269 43095 44327 43101
rect 44269 43092 44281 43095
rect 44232 43064 44281 43092
rect 44232 43052 44238 43064
rect 44269 43061 44281 43064
rect 44315 43061 44327 43095
rect 44269 43055 44327 43061
rect 45370 43052 45376 43104
rect 45428 43092 45434 43104
rect 46293 43095 46351 43101
rect 46293 43092 46305 43095
rect 45428 43064 46305 43092
rect 45428 43052 45434 43064
rect 46293 43061 46305 43064
rect 46339 43061 46351 43095
rect 46293 43055 46351 43061
rect 48130 43052 48136 43104
rect 48188 43092 48194 43104
rect 48225 43095 48283 43101
rect 48225 43092 48237 43095
rect 48188 43064 48237 43092
rect 48188 43052 48194 43064
rect 48225 43061 48237 43064
rect 48271 43092 48283 43095
rect 51046 43092 51074 43132
rect 53006 43120 53012 43132
rect 53064 43120 53070 43172
rect 52730 43092 52736 43104
rect 48271 43064 51074 43092
rect 52691 43064 52736 43092
rect 48271 43061 48283 43064
rect 48225 43055 48283 43061
rect 52730 43052 52736 43064
rect 52788 43052 52794 43104
rect 1104 43002 58880 43024
rect 1104 42950 4214 43002
rect 4266 42950 4278 43002
rect 4330 42950 4342 43002
rect 4394 42950 4406 43002
rect 4458 42950 4470 43002
rect 4522 42950 34934 43002
rect 34986 42950 34998 43002
rect 35050 42950 35062 43002
rect 35114 42950 35126 43002
rect 35178 42950 35190 43002
rect 35242 42950 58880 43002
rect 1104 42928 58880 42950
rect 38013 42891 38071 42897
rect 38013 42857 38025 42891
rect 38059 42888 38071 42891
rect 38286 42888 38292 42900
rect 38059 42860 38292 42888
rect 38059 42857 38071 42860
rect 38013 42851 38071 42857
rect 38286 42848 38292 42860
rect 38344 42848 38350 42900
rect 40037 42891 40095 42897
rect 40037 42857 40049 42891
rect 40083 42888 40095 42891
rect 40494 42888 40500 42900
rect 40083 42860 40500 42888
rect 40083 42857 40095 42860
rect 40037 42851 40095 42857
rect 40494 42848 40500 42860
rect 40552 42848 40558 42900
rect 45370 42888 45376 42900
rect 45331 42860 45376 42888
rect 45370 42848 45376 42860
rect 45428 42848 45434 42900
rect 49326 42848 49332 42900
rect 49384 42888 49390 42900
rect 49605 42891 49663 42897
rect 49605 42888 49617 42891
rect 49384 42860 49617 42888
rect 49384 42848 49390 42860
rect 49605 42857 49617 42860
rect 49651 42857 49663 42891
rect 49605 42851 49663 42857
rect 44453 42823 44511 42829
rect 44453 42789 44465 42823
rect 44499 42789 44511 42823
rect 47026 42820 47032 42832
rect 44453 42783 44511 42789
rect 45664 42792 47032 42820
rect 38654 42712 38660 42764
rect 38712 42752 38718 42764
rect 41371 42755 41429 42761
rect 41371 42752 41383 42755
rect 38712 42724 41383 42752
rect 38712 42712 38718 42724
rect 41371 42721 41383 42724
rect 41417 42721 41429 42755
rect 41371 42715 41429 42721
rect 41506 42712 41512 42764
rect 41564 42752 41570 42764
rect 41877 42755 41935 42761
rect 41877 42752 41889 42755
rect 41564 42724 41889 42752
rect 41564 42712 41570 42724
rect 41877 42721 41889 42724
rect 41923 42721 41935 42755
rect 44468 42752 44496 42783
rect 45281 42755 45339 42761
rect 45281 42752 45293 42755
rect 44468 42724 45293 42752
rect 41877 42715 41935 42721
rect 45281 42721 45293 42724
rect 45327 42752 45339 42755
rect 45554 42752 45560 42764
rect 45327 42724 45560 42752
rect 45327 42721 45339 42724
rect 45281 42715 45339 42721
rect 45554 42712 45560 42724
rect 45612 42712 45618 42764
rect 3973 42687 4031 42693
rect 3973 42653 3985 42687
rect 4019 42684 4031 42687
rect 9582 42684 9588 42696
rect 4019 42656 9588 42684
rect 4019 42653 4031 42656
rect 3973 42647 4031 42653
rect 9582 42644 9588 42656
rect 9640 42644 9646 42696
rect 36906 42693 36912 42696
rect 36633 42687 36691 42693
rect 36633 42653 36645 42687
rect 36679 42653 36691 42687
rect 36900 42684 36912 42693
rect 36867 42656 36912 42684
rect 36633 42647 36691 42653
rect 36900 42647 36912 42656
rect 36648 42616 36676 42647
rect 36906 42644 36912 42647
rect 36964 42644 36970 42696
rect 41141 42687 41199 42693
rect 41141 42653 41153 42687
rect 41187 42684 41199 42687
rect 41187 42656 43024 42684
rect 41187 42653 41199 42656
rect 41141 42647 41199 42653
rect 37274 42616 37280 42628
rect 36648 42588 37280 42616
rect 37274 42576 37280 42588
rect 37332 42576 37338 42628
rect 3881 42551 3939 42557
rect 3881 42517 3893 42551
rect 3927 42548 3939 42551
rect 3970 42548 3976 42560
rect 3927 42520 3976 42548
rect 3927 42517 3939 42520
rect 3881 42511 3939 42517
rect 3970 42508 3976 42520
rect 4028 42508 4034 42560
rect 41230 42508 41236 42560
rect 41288 42548 41294 42560
rect 41410 42551 41468 42557
rect 41410 42548 41422 42551
rect 41288 42520 41422 42548
rect 41288 42508 41294 42520
rect 41410 42517 41422 42520
rect 41456 42517 41468 42551
rect 42996 42548 43024 42656
rect 43070 42644 43076 42696
rect 43128 42684 43134 42696
rect 45373 42687 45431 42693
rect 43128 42656 43173 42684
rect 43128 42644 43134 42656
rect 45373 42653 45385 42687
rect 45419 42684 45431 42687
rect 45664 42684 45692 42792
rect 47026 42780 47032 42792
rect 47084 42780 47090 42832
rect 46014 42712 46020 42764
rect 46072 42761 46078 42764
rect 46072 42755 46094 42761
rect 46082 42721 46094 42755
rect 48222 42752 48228 42764
rect 48186 42724 48228 42752
rect 46072 42715 46094 42721
rect 46072 42712 46078 42715
rect 48222 42712 48228 42724
rect 48280 42712 48286 42764
rect 49418 42752 49424 42764
rect 48332 42724 49424 42752
rect 45830 42684 45836 42696
rect 45419 42656 45692 42684
rect 45791 42656 45836 42684
rect 45419 42653 45431 42656
rect 45373 42647 45431 42653
rect 45830 42644 45836 42656
rect 45888 42644 45894 42696
rect 45922 42644 45928 42696
rect 45980 42684 45986 42696
rect 47762 42684 47768 42696
rect 45980 42656 46025 42684
rect 47723 42656 47768 42684
rect 45980 42644 45986 42656
rect 47762 42644 47768 42656
rect 47820 42644 47826 42696
rect 48088 42687 48146 42693
rect 48088 42653 48100 42687
rect 48134 42684 48146 42687
rect 48332 42684 48360 42724
rect 49418 42712 49424 42724
rect 49476 42712 49482 42764
rect 48498 42684 48504 42696
rect 48134 42656 48360 42684
rect 48459 42656 48504 42684
rect 48134 42653 48146 42656
rect 48088 42647 48146 42653
rect 48498 42644 48504 42656
rect 48556 42644 48562 42696
rect 49620 42684 49648 42851
rect 50062 42848 50068 42900
rect 50120 42888 50126 42900
rect 50120 42860 51028 42888
rect 50120 42848 50126 42860
rect 50154 42712 50160 42764
rect 50212 42752 50218 42764
rect 50341 42755 50399 42761
rect 50341 42752 50353 42755
rect 50212 42724 50353 42752
rect 50212 42712 50218 42724
rect 50341 42721 50353 42724
rect 50387 42721 50399 42755
rect 51000 42752 51028 42860
rect 51813 42755 51871 42761
rect 51813 42752 51825 42755
rect 51000 42724 51825 42752
rect 50341 42715 50399 42721
rect 51813 42721 51825 42724
rect 51859 42721 51871 42755
rect 51813 42715 51871 42721
rect 52319 42755 52377 42761
rect 52319 42721 52331 42755
rect 52365 42752 52377 42755
rect 52638 42752 52644 42764
rect 52365 42724 52644 42752
rect 52365 42721 52377 42724
rect 52319 42715 52377 42721
rect 52638 42712 52644 42724
rect 52696 42712 52702 42764
rect 50617 42687 50675 42693
rect 50617 42684 50629 42687
rect 49620 42656 50629 42684
rect 50617 42653 50629 42656
rect 50663 42653 50675 42687
rect 52454 42684 52460 42696
rect 50617 42647 50675 42653
rect 51920 42656 52460 42684
rect 43340 42619 43398 42625
rect 43340 42585 43352 42619
rect 43386 42616 43398 42619
rect 43990 42616 43996 42628
rect 43386 42588 43996 42616
rect 43386 42585 43398 42588
rect 43340 42579 43398 42585
rect 43990 42576 43996 42588
rect 44048 42576 44054 42628
rect 44928 42588 46060 42616
rect 44928 42548 44956 42588
rect 42996 42520 44956 42548
rect 45005 42551 45063 42557
rect 41410 42511 41468 42517
rect 45005 42517 45017 42551
rect 45051 42548 45063 42551
rect 45554 42548 45560 42560
rect 45051 42520 45560 42548
rect 45051 42517 45063 42520
rect 45005 42511 45063 42517
rect 45554 42508 45560 42520
rect 45612 42508 45618 42560
rect 46032 42548 46060 42588
rect 46106 42576 46112 42628
rect 46164 42616 46170 42628
rect 46164 42588 46209 42616
rect 46164 42576 46170 42588
rect 48130 42548 48136 42560
rect 46032 42520 48136 42548
rect 48130 42508 48136 42520
rect 48188 42508 48194 42560
rect 51353 42551 51411 42557
rect 51353 42517 51365 42551
rect 51399 42548 51411 42551
rect 51920 42548 51948 42656
rect 52454 42644 52460 42656
rect 52512 42644 52518 42696
rect 52546 42644 52552 42696
rect 52604 42684 52610 42696
rect 52604 42656 52649 42684
rect 52604 42644 52610 42656
rect 56318 42644 56324 42696
rect 56376 42684 56382 42696
rect 57241 42687 57299 42693
rect 57241 42684 57253 42687
rect 56376 42656 57253 42684
rect 56376 42644 56382 42656
rect 57241 42653 57253 42656
rect 57287 42653 57299 42687
rect 57241 42647 57299 42653
rect 57054 42616 57060 42628
rect 53208 42588 57060 42616
rect 51399 42520 51948 42548
rect 51399 42517 51411 42520
rect 51353 42511 51411 42517
rect 52086 42508 52092 42560
rect 52144 42548 52150 42560
rect 52279 42551 52337 42557
rect 52279 42548 52291 42551
rect 52144 42520 52291 42548
rect 52144 42508 52150 42520
rect 52279 42517 52291 42520
rect 52325 42548 52337 42551
rect 53208 42548 53236 42588
rect 57054 42576 57060 42588
rect 57112 42576 57118 42628
rect 53650 42548 53656 42560
rect 52325 42520 53236 42548
rect 53611 42520 53656 42548
rect 52325 42517 52337 42520
rect 52279 42511 52337 42517
rect 53650 42508 53656 42520
rect 53708 42508 53714 42560
rect 1104 42458 58880 42480
rect 1104 42406 19574 42458
rect 19626 42406 19638 42458
rect 19690 42406 19702 42458
rect 19754 42406 19766 42458
rect 19818 42406 19830 42458
rect 19882 42406 50294 42458
rect 50346 42406 50358 42458
rect 50410 42406 50422 42458
rect 50474 42406 50486 42458
rect 50538 42406 50550 42458
rect 50602 42406 58880 42458
rect 1104 42384 58880 42406
rect 44174 42344 44180 42356
rect 44135 42316 44180 42344
rect 44174 42304 44180 42316
rect 44232 42304 44238 42356
rect 45462 42344 45468 42356
rect 44836 42316 45468 42344
rect 3970 42276 3976 42288
rect 3931 42248 3976 42276
rect 3970 42236 3976 42248
rect 4028 42236 4034 42288
rect 44836 42285 44864 42316
rect 45462 42304 45468 42316
rect 45520 42344 45526 42356
rect 46106 42344 46112 42356
rect 45520 42316 46112 42344
rect 45520 42304 45526 42316
rect 46106 42304 46112 42316
rect 46164 42304 46170 42356
rect 46937 42347 46995 42353
rect 46937 42313 46949 42347
rect 46983 42344 46995 42347
rect 47026 42344 47032 42356
rect 46983 42316 47032 42344
rect 46983 42313 46995 42316
rect 46937 42307 46995 42313
rect 47026 42304 47032 42316
rect 47084 42304 47090 42356
rect 48409 42347 48467 42353
rect 48409 42313 48421 42347
rect 48455 42344 48467 42347
rect 48498 42344 48504 42356
rect 48455 42316 48504 42344
rect 48455 42313 48467 42316
rect 48409 42307 48467 42313
rect 48498 42304 48504 42316
rect 48556 42344 48562 42356
rect 48556 42316 48912 42344
rect 48556 42304 48562 42316
rect 43993 42279 44051 42285
rect 43993 42245 44005 42279
rect 44039 42276 44051 42279
rect 44821 42279 44879 42285
rect 44821 42276 44833 42279
rect 44039 42248 44833 42276
rect 44039 42245 44051 42248
rect 43993 42239 44051 42245
rect 44821 42245 44833 42248
rect 44867 42245 44879 42279
rect 44821 42239 44879 42245
rect 45005 42279 45063 42285
rect 45005 42245 45017 42279
rect 45051 42276 45063 42279
rect 45554 42276 45560 42288
rect 45051 42248 45560 42276
rect 45051 42245 45063 42248
rect 45005 42239 45063 42245
rect 45554 42236 45560 42248
rect 45612 42236 45618 42288
rect 4154 42168 4160 42220
rect 4212 42208 4218 42220
rect 4212 42180 4257 42208
rect 4212 42168 4218 42180
rect 44266 42168 44272 42220
rect 44324 42208 44330 42220
rect 44324 42180 44369 42208
rect 44324 42168 44330 42180
rect 45094 42168 45100 42220
rect 45152 42208 45158 42220
rect 45813 42211 45871 42217
rect 45813 42208 45825 42211
rect 45152 42180 45197 42208
rect 45296 42180 45825 42208
rect 45152 42168 45158 42180
rect 2774 42140 2780 42152
rect 2735 42112 2780 42140
rect 2774 42100 2780 42112
rect 2832 42100 2838 42152
rect 9582 42032 9588 42084
rect 9640 42072 9646 42084
rect 33594 42072 33600 42084
rect 9640 42044 33600 42072
rect 9640 42032 9646 42044
rect 33594 42032 33600 42044
rect 33652 42032 33658 42084
rect 43990 42072 43996 42084
rect 43951 42044 43996 42072
rect 43990 42032 43996 42044
rect 44048 42032 44054 42084
rect 44821 42075 44879 42081
rect 44821 42041 44833 42075
rect 44867 42072 44879 42075
rect 45296 42072 45324 42180
rect 45813 42177 45825 42180
rect 45859 42177 45871 42211
rect 48884 42208 48912 42316
rect 49418 42304 49424 42356
rect 49476 42344 49482 42356
rect 49782 42347 49840 42353
rect 49782 42344 49794 42347
rect 49476 42316 49794 42344
rect 49476 42304 49482 42316
rect 49782 42313 49794 42316
rect 49828 42344 49840 42347
rect 51994 42344 52000 42356
rect 49828 42316 52000 42344
rect 49828 42313 49840 42316
rect 49782 42307 49840 42313
rect 51994 42304 52000 42316
rect 52052 42304 52058 42356
rect 52089 42347 52147 42353
rect 52089 42313 52101 42347
rect 52135 42344 52147 42347
rect 52822 42344 52828 42356
rect 52135 42316 52828 42344
rect 52135 42313 52147 42316
rect 52089 42307 52147 42313
rect 52822 42304 52828 42316
rect 52880 42304 52886 42356
rect 52914 42304 52920 42356
rect 52972 42344 52978 42356
rect 53745 42347 53803 42353
rect 53745 42344 53757 42347
rect 52972 42316 53757 42344
rect 52972 42304 52978 42316
rect 53745 42313 53757 42316
rect 53791 42313 53803 42347
rect 53745 42307 53803 42313
rect 51353 42211 51411 42217
rect 51353 42208 51365 42211
rect 48884 42180 51365 42208
rect 45813 42171 45871 42177
rect 51353 42177 51365 42180
rect 51399 42177 51411 42211
rect 53006 42208 53012 42220
rect 52967 42180 53012 42208
rect 51353 42171 51411 42177
rect 53006 42168 53012 42180
rect 53064 42168 53070 42220
rect 56870 42208 56876 42220
rect 56831 42180 56876 42208
rect 56870 42168 56876 42180
rect 56928 42168 56934 42220
rect 45557 42143 45615 42149
rect 45557 42109 45569 42143
rect 45603 42109 45615 42143
rect 49510 42140 49516 42152
rect 49471 42112 49516 42140
rect 45557 42103 45615 42109
rect 44867 42044 45324 42072
rect 44867 42041 44879 42044
rect 44821 42035 44879 42041
rect 43070 41964 43076 42016
rect 43128 42004 43134 42016
rect 45572 42004 45600 42103
rect 49510 42100 49516 42112
rect 49568 42100 49574 42152
rect 49694 42100 49700 42152
rect 49752 42140 49758 42152
rect 49786 42143 49844 42149
rect 49786 42140 49798 42143
rect 49752 42112 49798 42140
rect 49752 42100 49758 42112
rect 49786 42109 49798 42112
rect 49832 42109 49844 42143
rect 49786 42103 49844 42109
rect 50062 42100 50068 42152
rect 50120 42140 50126 42152
rect 50249 42143 50307 42149
rect 50249 42140 50261 42143
rect 50120 42112 50261 42140
rect 50120 42100 50126 42112
rect 50249 42109 50261 42112
rect 50295 42109 50307 42143
rect 50249 42103 50307 42109
rect 50338 42100 50344 42152
rect 50396 42140 50402 42152
rect 51074 42140 51080 42152
rect 50396 42112 51080 42140
rect 50396 42100 50402 42112
rect 51074 42100 51080 42112
rect 51132 42100 51138 42152
rect 51718 42100 51724 42152
rect 51776 42140 51782 42152
rect 52733 42143 52791 42149
rect 52733 42140 52745 42143
rect 51776 42112 52745 42140
rect 51776 42100 51782 42112
rect 52733 42109 52745 42112
rect 52779 42109 52791 42143
rect 52733 42103 52791 42109
rect 45738 42004 45744 42016
rect 43128 41976 45744 42004
rect 43128 41964 43134 41976
rect 45738 41964 45744 41976
rect 45796 41964 45802 42016
rect 47762 41964 47768 42016
rect 47820 42004 47826 42016
rect 50062 42004 50068 42016
rect 47820 41976 50068 42004
rect 47820 41964 47826 41976
rect 50062 41964 50068 41976
rect 50120 41964 50126 42016
rect 56502 41964 56508 42016
rect 56560 42004 56566 42016
rect 56781 42007 56839 42013
rect 56781 42004 56793 42007
rect 56560 41976 56793 42004
rect 56560 41964 56566 41976
rect 56781 41973 56793 41976
rect 56827 41973 56839 42007
rect 56781 41967 56839 41973
rect 1104 41914 58880 41936
rect 1104 41862 4214 41914
rect 4266 41862 4278 41914
rect 4330 41862 4342 41914
rect 4394 41862 4406 41914
rect 4458 41862 4470 41914
rect 4522 41862 34934 41914
rect 34986 41862 34998 41914
rect 35050 41862 35062 41914
rect 35114 41862 35126 41914
rect 35178 41862 35190 41914
rect 35242 41862 58880 41914
rect 1104 41840 58880 41862
rect 45094 41800 45100 41812
rect 45055 41772 45100 41800
rect 45094 41760 45100 41772
rect 45152 41760 45158 41812
rect 46934 41760 46940 41812
rect 46992 41800 46998 41812
rect 47118 41800 47124 41812
rect 46992 41772 47124 41800
rect 46992 41760 46998 41772
rect 47118 41760 47124 41772
rect 47176 41760 47182 41812
rect 52730 41800 52736 41812
rect 52691 41772 52736 41800
rect 52730 41760 52736 41772
rect 52788 41760 52794 41812
rect 45738 41664 45744 41676
rect 45699 41636 45744 41664
rect 45738 41624 45744 41636
rect 45796 41624 45802 41676
rect 51074 41624 51080 41676
rect 51132 41664 51138 41676
rect 51718 41664 51724 41676
rect 51132 41636 51724 41664
rect 51132 41624 51138 41636
rect 51718 41624 51724 41636
rect 51776 41624 51782 41676
rect 56318 41664 56324 41676
rect 56279 41636 56324 41664
rect 56318 41624 56324 41636
rect 56376 41624 56382 41676
rect 56502 41664 56508 41676
rect 56463 41636 56508 41664
rect 56502 41624 56508 41636
rect 56560 41624 56566 41676
rect 58158 41664 58164 41676
rect 58119 41636 58164 41664
rect 58158 41624 58164 41636
rect 58216 41624 58222 41676
rect 44174 41556 44180 41608
rect 44232 41596 44238 41608
rect 46014 41605 46020 41608
rect 45005 41599 45063 41605
rect 45005 41596 45017 41599
rect 44232 41568 45017 41596
rect 44232 41556 44238 41568
rect 45005 41565 45017 41568
rect 45051 41565 45063 41599
rect 45005 41559 45063 41565
rect 45189 41599 45247 41605
rect 45189 41565 45201 41599
rect 45235 41565 45247 41599
rect 46008 41596 46020 41605
rect 45975 41568 46020 41596
rect 45189 41559 45247 41565
rect 46008 41559 46020 41568
rect 45204 41528 45232 41559
rect 46014 41556 46020 41559
rect 46072 41556 46078 41608
rect 51997 41599 52055 41605
rect 51997 41565 52009 41599
rect 52043 41596 52055 41599
rect 53650 41596 53656 41608
rect 52043 41568 53656 41596
rect 52043 41565 52055 41568
rect 51997 41559 52055 41565
rect 47026 41528 47032 41540
rect 45204 41500 47032 41528
rect 47026 41488 47032 41500
rect 47084 41488 47090 41540
rect 49510 41488 49516 41540
rect 49568 41528 49574 41540
rect 52012 41528 52040 41559
rect 53650 41556 53656 41568
rect 53708 41556 53714 41608
rect 49568 41500 52040 41528
rect 49568 41488 49574 41500
rect 1104 41370 58880 41392
rect 1104 41318 19574 41370
rect 19626 41318 19638 41370
rect 19690 41318 19702 41370
rect 19754 41318 19766 41370
rect 19818 41318 19830 41370
rect 19882 41318 50294 41370
rect 50346 41318 50358 41370
rect 50410 41318 50422 41370
rect 50474 41318 50486 41370
rect 50538 41318 50550 41370
rect 50602 41318 58880 41370
rect 1104 41296 58880 41318
rect 45741 41259 45799 41265
rect 45741 41225 45753 41259
rect 45787 41256 45799 41259
rect 45830 41256 45836 41268
rect 45787 41228 45836 41256
rect 45787 41225 45799 41228
rect 45741 41219 45799 41225
rect 45830 41216 45836 41228
rect 45888 41216 45894 41268
rect 45554 41080 45560 41132
rect 45612 41120 45618 41132
rect 45741 41123 45799 41129
rect 45612 41092 45657 41120
rect 45612 41080 45618 41092
rect 45741 41089 45753 41123
rect 45787 41120 45799 41123
rect 47118 41120 47124 41132
rect 45787 41092 47124 41120
rect 45787 41089 45799 41092
rect 45741 41083 45799 41089
rect 47118 41080 47124 41092
rect 47176 41080 47182 41132
rect 1104 40826 58880 40848
rect 1104 40774 4214 40826
rect 4266 40774 4278 40826
rect 4330 40774 4342 40826
rect 4394 40774 4406 40826
rect 4458 40774 4470 40826
rect 4522 40774 34934 40826
rect 34986 40774 34998 40826
rect 35050 40774 35062 40826
rect 35114 40774 35126 40826
rect 35178 40774 35190 40826
rect 35242 40774 58880 40826
rect 1104 40752 58880 40774
rect 1104 40282 58880 40304
rect 1104 40230 19574 40282
rect 19626 40230 19638 40282
rect 19690 40230 19702 40282
rect 19754 40230 19766 40282
rect 19818 40230 19830 40282
rect 19882 40230 50294 40282
rect 50346 40230 50358 40282
rect 50410 40230 50422 40282
rect 50474 40230 50486 40282
rect 50538 40230 50550 40282
rect 50602 40230 58880 40282
rect 1104 40208 58880 40230
rect 1104 39738 58880 39760
rect 1104 39686 4214 39738
rect 4266 39686 4278 39738
rect 4330 39686 4342 39738
rect 4394 39686 4406 39738
rect 4458 39686 4470 39738
rect 4522 39686 34934 39738
rect 34986 39686 34998 39738
rect 35050 39686 35062 39738
rect 35114 39686 35126 39738
rect 35178 39686 35190 39738
rect 35242 39686 58880 39738
rect 1104 39664 58880 39686
rect 1104 39194 58880 39216
rect 1104 39142 19574 39194
rect 19626 39142 19638 39194
rect 19690 39142 19702 39194
rect 19754 39142 19766 39194
rect 19818 39142 19830 39194
rect 19882 39142 50294 39194
rect 50346 39142 50358 39194
rect 50410 39142 50422 39194
rect 50474 39142 50486 39194
rect 50538 39142 50550 39194
rect 50602 39142 58880 39194
rect 1104 39120 58880 39142
rect 1104 38650 58880 38672
rect 1104 38598 4214 38650
rect 4266 38598 4278 38650
rect 4330 38598 4342 38650
rect 4394 38598 4406 38650
rect 4458 38598 4470 38650
rect 4522 38598 34934 38650
rect 34986 38598 34998 38650
rect 35050 38598 35062 38650
rect 35114 38598 35126 38650
rect 35178 38598 35190 38650
rect 35242 38598 58880 38650
rect 1104 38576 58880 38598
rect 1104 38106 58880 38128
rect 1104 38054 19574 38106
rect 19626 38054 19638 38106
rect 19690 38054 19702 38106
rect 19754 38054 19766 38106
rect 19818 38054 19830 38106
rect 19882 38054 50294 38106
rect 50346 38054 50358 38106
rect 50410 38054 50422 38106
rect 50474 38054 50486 38106
rect 50538 38054 50550 38106
rect 50602 38054 58880 38106
rect 1104 38032 58880 38054
rect 1104 37562 58880 37584
rect 1104 37510 4214 37562
rect 4266 37510 4278 37562
rect 4330 37510 4342 37562
rect 4394 37510 4406 37562
rect 4458 37510 4470 37562
rect 4522 37510 34934 37562
rect 34986 37510 34998 37562
rect 35050 37510 35062 37562
rect 35114 37510 35126 37562
rect 35178 37510 35190 37562
rect 35242 37510 58880 37562
rect 1104 37488 58880 37510
rect 1104 37018 58880 37040
rect 1104 36966 19574 37018
rect 19626 36966 19638 37018
rect 19690 36966 19702 37018
rect 19754 36966 19766 37018
rect 19818 36966 19830 37018
rect 19882 36966 50294 37018
rect 50346 36966 50358 37018
rect 50410 36966 50422 37018
rect 50474 36966 50486 37018
rect 50538 36966 50550 37018
rect 50602 36966 58880 37018
rect 1104 36944 58880 36966
rect 1104 36474 58880 36496
rect 1104 36422 4214 36474
rect 4266 36422 4278 36474
rect 4330 36422 4342 36474
rect 4394 36422 4406 36474
rect 4458 36422 4470 36474
rect 4522 36422 34934 36474
rect 34986 36422 34998 36474
rect 35050 36422 35062 36474
rect 35114 36422 35126 36474
rect 35178 36422 35190 36474
rect 35242 36422 58880 36474
rect 1104 36400 58880 36422
rect 1104 35930 58880 35952
rect 1104 35878 19574 35930
rect 19626 35878 19638 35930
rect 19690 35878 19702 35930
rect 19754 35878 19766 35930
rect 19818 35878 19830 35930
rect 19882 35878 50294 35930
rect 50346 35878 50358 35930
rect 50410 35878 50422 35930
rect 50474 35878 50486 35930
rect 50538 35878 50550 35930
rect 50602 35878 58880 35930
rect 1104 35856 58880 35878
rect 1104 35386 58880 35408
rect 1104 35334 4214 35386
rect 4266 35334 4278 35386
rect 4330 35334 4342 35386
rect 4394 35334 4406 35386
rect 4458 35334 4470 35386
rect 4522 35334 34934 35386
rect 34986 35334 34998 35386
rect 35050 35334 35062 35386
rect 35114 35334 35126 35386
rect 35178 35334 35190 35386
rect 35242 35334 58880 35386
rect 1104 35312 58880 35334
rect 2406 35068 2412 35080
rect 2367 35040 2412 35068
rect 2406 35028 2412 35040
rect 2464 35028 2470 35080
rect 3973 35071 4031 35077
rect 3973 35037 3985 35071
rect 4019 35068 4031 35071
rect 4614 35068 4620 35080
rect 4019 35040 4620 35068
rect 4019 35037 4031 35040
rect 3973 35031 4031 35037
rect 4614 35028 4620 35040
rect 4672 35068 4678 35080
rect 9030 35068 9036 35080
rect 4672 35040 9036 35068
rect 4672 35028 4678 35040
rect 9030 35028 9036 35040
rect 9088 35028 9094 35080
rect 3786 34892 3792 34944
rect 3844 34932 3850 34944
rect 3881 34935 3939 34941
rect 3881 34932 3893 34935
rect 3844 34904 3893 34932
rect 3844 34892 3850 34904
rect 3881 34901 3893 34904
rect 3927 34901 3939 34935
rect 3881 34895 3939 34901
rect 1104 34842 58880 34864
rect 1104 34790 19574 34842
rect 19626 34790 19638 34842
rect 19690 34790 19702 34842
rect 19754 34790 19766 34842
rect 19818 34790 19830 34842
rect 19882 34790 50294 34842
rect 50346 34790 50358 34842
rect 50410 34790 50422 34842
rect 50474 34790 50486 34842
rect 50538 34790 50550 34842
rect 50602 34790 58880 34842
rect 1104 34768 58880 34790
rect 2130 34660 2136 34672
rect 2091 34632 2136 34660
rect 2130 34620 2136 34632
rect 2188 34620 2194 34672
rect 3786 34660 3792 34672
rect 3747 34632 3792 34660
rect 3786 34620 3792 34632
rect 3844 34620 3850 34672
rect 2406 34484 2412 34536
rect 2464 34524 2470 34536
rect 3973 34527 4031 34533
rect 3973 34524 3985 34527
rect 2464 34496 3985 34524
rect 2464 34484 2470 34496
rect 3973 34493 3985 34496
rect 4019 34493 4031 34527
rect 3973 34487 4031 34493
rect 1104 34298 58880 34320
rect 1104 34246 4214 34298
rect 4266 34246 4278 34298
rect 4330 34246 4342 34298
rect 4394 34246 4406 34298
rect 4458 34246 4470 34298
rect 4522 34246 34934 34298
rect 34986 34246 34998 34298
rect 35050 34246 35062 34298
rect 35114 34246 35126 34298
rect 35178 34246 35190 34298
rect 35242 34246 58880 34298
rect 1104 34224 58880 34246
rect 1104 33754 58880 33776
rect 1104 33702 19574 33754
rect 19626 33702 19638 33754
rect 19690 33702 19702 33754
rect 19754 33702 19766 33754
rect 19818 33702 19830 33754
rect 19882 33702 50294 33754
rect 50346 33702 50358 33754
rect 50410 33702 50422 33754
rect 50474 33702 50486 33754
rect 50538 33702 50550 33754
rect 50602 33702 58880 33754
rect 1104 33680 58880 33702
rect 1104 33210 58880 33232
rect 1104 33158 4214 33210
rect 4266 33158 4278 33210
rect 4330 33158 4342 33210
rect 4394 33158 4406 33210
rect 4458 33158 4470 33210
rect 4522 33158 34934 33210
rect 34986 33158 34998 33210
rect 35050 33158 35062 33210
rect 35114 33158 35126 33210
rect 35178 33158 35190 33210
rect 35242 33158 58880 33210
rect 1104 33136 58880 33158
rect 1104 32666 58880 32688
rect 1104 32614 19574 32666
rect 19626 32614 19638 32666
rect 19690 32614 19702 32666
rect 19754 32614 19766 32666
rect 19818 32614 19830 32666
rect 19882 32614 50294 32666
rect 50346 32614 50358 32666
rect 50410 32614 50422 32666
rect 50474 32614 50486 32666
rect 50538 32614 50550 32666
rect 50602 32614 58880 32666
rect 1104 32592 58880 32614
rect 1104 32122 58880 32144
rect 1104 32070 4214 32122
rect 4266 32070 4278 32122
rect 4330 32070 4342 32122
rect 4394 32070 4406 32122
rect 4458 32070 4470 32122
rect 4522 32070 34934 32122
rect 34986 32070 34998 32122
rect 35050 32070 35062 32122
rect 35114 32070 35126 32122
rect 35178 32070 35190 32122
rect 35242 32070 58880 32122
rect 1104 32048 58880 32070
rect 57054 31872 57060 31884
rect 57015 31844 57060 31872
rect 57054 31832 57060 31844
rect 57112 31832 57118 31884
rect 58158 31804 58164 31816
rect 58119 31776 58164 31804
rect 58158 31764 58164 31776
rect 58216 31764 58222 31816
rect 1104 31578 58880 31600
rect 1104 31526 19574 31578
rect 19626 31526 19638 31578
rect 19690 31526 19702 31578
rect 19754 31526 19766 31578
rect 19818 31526 19830 31578
rect 19882 31526 50294 31578
rect 50346 31526 50358 31578
rect 50410 31526 50422 31578
rect 50474 31526 50486 31578
rect 50538 31526 50550 31578
rect 50602 31526 58880 31578
rect 1104 31504 58880 31526
rect 1104 31034 58880 31056
rect 1104 30982 4214 31034
rect 4266 30982 4278 31034
rect 4330 30982 4342 31034
rect 4394 30982 4406 31034
rect 4458 30982 4470 31034
rect 4522 30982 34934 31034
rect 34986 30982 34998 31034
rect 35050 30982 35062 31034
rect 35114 30982 35126 31034
rect 35178 30982 35190 31034
rect 35242 30982 58880 31034
rect 1104 30960 58880 30982
rect 1104 30490 58880 30512
rect 1104 30438 19574 30490
rect 19626 30438 19638 30490
rect 19690 30438 19702 30490
rect 19754 30438 19766 30490
rect 19818 30438 19830 30490
rect 19882 30438 50294 30490
rect 50346 30438 50358 30490
rect 50410 30438 50422 30490
rect 50474 30438 50486 30490
rect 50538 30438 50550 30490
rect 50602 30438 58880 30490
rect 1104 30416 58880 30438
rect 1104 29946 58880 29968
rect 1104 29894 4214 29946
rect 4266 29894 4278 29946
rect 4330 29894 4342 29946
rect 4394 29894 4406 29946
rect 4458 29894 4470 29946
rect 4522 29894 34934 29946
rect 34986 29894 34998 29946
rect 35050 29894 35062 29946
rect 35114 29894 35126 29946
rect 35178 29894 35190 29946
rect 35242 29894 58880 29946
rect 1104 29872 58880 29894
rect 1104 29402 58880 29424
rect 1104 29350 19574 29402
rect 19626 29350 19638 29402
rect 19690 29350 19702 29402
rect 19754 29350 19766 29402
rect 19818 29350 19830 29402
rect 19882 29350 50294 29402
rect 50346 29350 50358 29402
rect 50410 29350 50422 29402
rect 50474 29350 50486 29402
rect 50538 29350 50550 29402
rect 50602 29350 58880 29402
rect 1104 29328 58880 29350
rect 56962 29152 56968 29164
rect 56923 29124 56968 29152
rect 56962 29112 56968 29124
rect 57020 29112 57026 29164
rect 57057 29019 57115 29025
rect 57057 28985 57069 29019
rect 57103 29016 57115 29019
rect 57974 29016 57980 29028
rect 57103 28988 57980 29016
rect 57103 28985 57115 28988
rect 57057 28979 57115 28985
rect 57974 28976 57980 28988
rect 58032 28976 58038 29028
rect 58069 28951 58127 28957
rect 58069 28917 58081 28951
rect 58115 28948 58127 28951
rect 58158 28948 58164 28960
rect 58115 28920 58164 28948
rect 58115 28917 58127 28920
rect 58069 28911 58127 28917
rect 58158 28908 58164 28920
rect 58216 28908 58222 28960
rect 1104 28858 58880 28880
rect 1104 28806 4214 28858
rect 4266 28806 4278 28858
rect 4330 28806 4342 28858
rect 4394 28806 4406 28858
rect 4458 28806 4470 28858
rect 4522 28806 34934 28858
rect 34986 28806 34998 28858
rect 35050 28806 35062 28858
rect 35114 28806 35126 28858
rect 35178 28806 35190 28858
rect 35242 28806 58880 28858
rect 1104 28784 58880 28806
rect 57698 28608 57704 28620
rect 57659 28580 57704 28608
rect 57698 28568 57704 28580
rect 57756 28568 57762 28620
rect 57974 28608 57980 28620
rect 57935 28580 57980 28608
rect 57974 28568 57980 28580
rect 58032 28568 58038 28620
rect 58158 28608 58164 28620
rect 58119 28580 58164 28608
rect 58158 28568 58164 28580
rect 58216 28568 58222 28620
rect 1104 28314 58880 28336
rect 1104 28262 19574 28314
rect 19626 28262 19638 28314
rect 19690 28262 19702 28314
rect 19754 28262 19766 28314
rect 19818 28262 19830 28314
rect 19882 28262 50294 28314
rect 50346 28262 50358 28314
rect 50410 28262 50422 28314
rect 50474 28262 50486 28314
rect 50538 28262 50550 28314
rect 50602 28262 58880 28314
rect 1104 28240 58880 28262
rect 1104 27770 58880 27792
rect 1104 27718 4214 27770
rect 4266 27718 4278 27770
rect 4330 27718 4342 27770
rect 4394 27718 4406 27770
rect 4458 27718 4470 27770
rect 4522 27718 34934 27770
rect 34986 27718 34998 27770
rect 35050 27718 35062 27770
rect 35114 27718 35126 27770
rect 35178 27718 35190 27770
rect 35242 27718 58880 27770
rect 1104 27696 58880 27718
rect 1104 27226 58880 27248
rect 1104 27174 19574 27226
rect 19626 27174 19638 27226
rect 19690 27174 19702 27226
rect 19754 27174 19766 27226
rect 19818 27174 19830 27226
rect 19882 27174 50294 27226
rect 50346 27174 50358 27226
rect 50410 27174 50422 27226
rect 50474 27174 50486 27226
rect 50538 27174 50550 27226
rect 50602 27174 58880 27226
rect 1104 27152 58880 27174
rect 1104 26682 58880 26704
rect 1104 26630 4214 26682
rect 4266 26630 4278 26682
rect 4330 26630 4342 26682
rect 4394 26630 4406 26682
rect 4458 26630 4470 26682
rect 4522 26630 34934 26682
rect 34986 26630 34998 26682
rect 35050 26630 35062 26682
rect 35114 26630 35126 26682
rect 35178 26630 35190 26682
rect 35242 26630 58880 26682
rect 1104 26608 58880 26630
rect 1104 26138 58880 26160
rect 1104 26086 19574 26138
rect 19626 26086 19638 26138
rect 19690 26086 19702 26138
rect 19754 26086 19766 26138
rect 19818 26086 19830 26138
rect 19882 26086 50294 26138
rect 50346 26086 50358 26138
rect 50410 26086 50422 26138
rect 50474 26086 50486 26138
rect 50538 26086 50550 26138
rect 50602 26086 58880 26138
rect 1104 26064 58880 26086
rect 8202 26024 8208 26036
rect 8163 25996 8208 26024
rect 8202 25984 8208 25996
rect 8260 25984 8266 26036
rect 8294 25888 8300 25900
rect 8255 25860 8300 25888
rect 8294 25848 8300 25860
rect 8352 25848 8358 25900
rect 1104 25594 58880 25616
rect 1104 25542 4214 25594
rect 4266 25542 4278 25594
rect 4330 25542 4342 25594
rect 4394 25542 4406 25594
rect 4458 25542 4470 25594
rect 4522 25542 34934 25594
rect 34986 25542 34998 25594
rect 35050 25542 35062 25594
rect 35114 25542 35126 25594
rect 35178 25542 35190 25594
rect 35242 25542 58880 25594
rect 1104 25520 58880 25542
rect 1104 25050 58880 25072
rect 1104 24998 19574 25050
rect 19626 24998 19638 25050
rect 19690 24998 19702 25050
rect 19754 24998 19766 25050
rect 19818 24998 19830 25050
rect 19882 24998 50294 25050
rect 50346 24998 50358 25050
rect 50410 24998 50422 25050
rect 50474 24998 50486 25050
rect 50538 24998 50550 25050
rect 50602 24998 58880 25050
rect 1104 24976 58880 24998
rect 8294 24760 8300 24812
rect 8352 24800 8358 24812
rect 8941 24803 8999 24809
rect 8941 24800 8953 24803
rect 8352 24772 8953 24800
rect 8352 24760 8358 24772
rect 8941 24769 8953 24772
rect 8987 24800 8999 24803
rect 55585 24803 55643 24809
rect 55585 24800 55597 24803
rect 8987 24772 55597 24800
rect 8987 24769 8999 24772
rect 8941 24763 8999 24769
rect 55585 24769 55597 24772
rect 55631 24800 55643 24803
rect 57054 24800 57060 24812
rect 55631 24772 57060 24800
rect 55631 24769 55643 24772
rect 55585 24763 55643 24769
rect 57054 24760 57060 24772
rect 57112 24760 57118 24812
rect 9582 24692 9588 24744
rect 9640 24732 9646 24744
rect 9953 24735 10011 24741
rect 9953 24732 9965 24735
rect 9640 24704 9965 24732
rect 9640 24692 9646 24704
rect 9953 24701 9965 24704
rect 9999 24732 10011 24735
rect 56226 24732 56232 24744
rect 9999 24704 45554 24732
rect 56187 24704 56232 24732
rect 9999 24701 10011 24704
rect 9953 24695 10011 24701
rect 45526 24664 45554 24704
rect 56226 24692 56232 24704
rect 56284 24692 56290 24744
rect 57790 24664 57796 24676
rect 45526 24636 57796 24664
rect 57790 24624 57796 24636
rect 57848 24624 57854 24676
rect 56502 24556 56508 24608
rect 56560 24596 56566 24608
rect 56965 24599 57023 24605
rect 56965 24596 56977 24599
rect 56560 24568 56977 24596
rect 56560 24556 56566 24568
rect 56965 24565 56977 24568
rect 57011 24565 57023 24599
rect 57882 24596 57888 24608
rect 57843 24568 57888 24596
rect 56965 24559 57023 24565
rect 57882 24556 57888 24568
rect 57940 24556 57946 24608
rect 1104 24506 58880 24528
rect 1104 24454 4214 24506
rect 4266 24454 4278 24506
rect 4330 24454 4342 24506
rect 4394 24454 4406 24506
rect 4458 24454 4470 24506
rect 4522 24454 34934 24506
rect 34986 24454 34998 24506
rect 35050 24454 35062 24506
rect 35114 24454 35126 24506
rect 35178 24454 35190 24506
rect 35242 24454 58880 24506
rect 1104 24432 58880 24454
rect 57882 24324 57888 24336
rect 56336 24296 57888 24324
rect 56336 24265 56364 24296
rect 57882 24284 57888 24296
rect 57940 24284 57946 24336
rect 56321 24259 56379 24265
rect 56321 24225 56333 24259
rect 56367 24225 56379 24259
rect 56502 24256 56508 24268
rect 56463 24228 56508 24256
rect 56321 24219 56379 24225
rect 56502 24216 56508 24228
rect 56560 24216 56566 24268
rect 58158 24256 58164 24268
rect 58119 24228 58164 24256
rect 58158 24216 58164 24228
rect 58216 24216 58222 24268
rect 1104 23962 58880 23984
rect 1104 23910 19574 23962
rect 19626 23910 19638 23962
rect 19690 23910 19702 23962
rect 19754 23910 19766 23962
rect 19818 23910 19830 23962
rect 19882 23910 50294 23962
rect 50346 23910 50358 23962
rect 50410 23910 50422 23962
rect 50474 23910 50486 23962
rect 50538 23910 50550 23962
rect 50602 23910 58880 23962
rect 1104 23888 58880 23910
rect 57054 23780 57060 23792
rect 57015 23752 57060 23780
rect 57054 23740 57060 23752
rect 57112 23740 57118 23792
rect 55585 23511 55643 23517
rect 55585 23477 55597 23511
rect 55631 23508 55643 23511
rect 55674 23508 55680 23520
rect 55631 23480 55680 23508
rect 55631 23477 55643 23480
rect 55585 23471 55643 23477
rect 55674 23468 55680 23480
rect 55732 23468 55738 23520
rect 1104 23418 58880 23440
rect 1104 23366 4214 23418
rect 4266 23366 4278 23418
rect 4330 23366 4342 23418
rect 4394 23366 4406 23418
rect 4458 23366 4470 23418
rect 4522 23366 34934 23418
rect 34986 23366 34998 23418
rect 35050 23366 35062 23418
rect 35114 23366 35126 23418
rect 35178 23366 35190 23418
rect 35242 23366 58880 23418
rect 1104 23344 58880 23366
rect 8205 23171 8263 23177
rect 8205 23137 8217 23171
rect 8251 23168 8263 23171
rect 8294 23168 8300 23180
rect 8251 23140 8300 23168
rect 8251 23137 8263 23140
rect 8205 23131 8263 23137
rect 8294 23128 8300 23140
rect 8352 23128 8358 23180
rect 7558 23060 7564 23112
rect 7616 23100 7622 23112
rect 7745 23103 7803 23109
rect 7745 23100 7757 23103
rect 7616 23072 7757 23100
rect 7616 23060 7622 23072
rect 7745 23069 7757 23072
rect 7791 23069 7803 23103
rect 7745 23063 7803 23069
rect 1104 22874 58880 22896
rect 1104 22822 19574 22874
rect 19626 22822 19638 22874
rect 19690 22822 19702 22874
rect 19754 22822 19766 22874
rect 19818 22822 19830 22874
rect 19882 22822 50294 22874
rect 50346 22822 50358 22874
rect 50410 22822 50422 22874
rect 50474 22822 50486 22874
rect 50538 22822 50550 22874
rect 50602 22822 58880 22874
rect 1104 22800 58880 22822
rect 7558 22624 7564 22636
rect 7519 22596 7564 22624
rect 7558 22584 7564 22596
rect 7616 22584 7622 22636
rect 8846 22420 8852 22432
rect 8807 22392 8852 22420
rect 8846 22380 8852 22392
rect 8904 22420 8910 22432
rect 56962 22420 56968 22432
rect 8904 22392 56968 22420
rect 8904 22380 8910 22392
rect 56962 22380 56968 22392
rect 57020 22380 57026 22432
rect 1104 22330 58880 22352
rect 1104 22278 4214 22330
rect 4266 22278 4278 22330
rect 4330 22278 4342 22330
rect 4394 22278 4406 22330
rect 4458 22278 4470 22330
rect 4522 22278 34934 22330
rect 34986 22278 34998 22330
rect 35050 22278 35062 22330
rect 35114 22278 35126 22330
rect 35178 22278 35190 22330
rect 35242 22278 58880 22330
rect 1104 22256 58880 22278
rect 1104 21786 58880 21808
rect 1104 21734 19574 21786
rect 19626 21734 19638 21786
rect 19690 21734 19702 21786
rect 19754 21734 19766 21786
rect 19818 21734 19830 21786
rect 19882 21734 50294 21786
rect 50346 21734 50358 21786
rect 50410 21734 50422 21786
rect 50474 21734 50486 21786
rect 50538 21734 50550 21786
rect 50602 21734 58880 21786
rect 1104 21712 58880 21734
rect 1104 21242 58880 21264
rect 1104 21190 4214 21242
rect 4266 21190 4278 21242
rect 4330 21190 4342 21242
rect 4394 21190 4406 21242
rect 4458 21190 4470 21242
rect 4522 21190 34934 21242
rect 34986 21190 34998 21242
rect 35050 21190 35062 21242
rect 35114 21190 35126 21242
rect 35178 21190 35190 21242
rect 35242 21190 58880 21242
rect 1104 21168 58880 21190
rect 1104 20698 58880 20720
rect 1104 20646 19574 20698
rect 19626 20646 19638 20698
rect 19690 20646 19702 20698
rect 19754 20646 19766 20698
rect 19818 20646 19830 20698
rect 19882 20646 50294 20698
rect 50346 20646 50358 20698
rect 50410 20646 50422 20698
rect 50474 20646 50486 20698
rect 50538 20646 50550 20698
rect 50602 20646 58880 20698
rect 1104 20624 58880 20646
rect 1104 20154 58880 20176
rect 1104 20102 4214 20154
rect 4266 20102 4278 20154
rect 4330 20102 4342 20154
rect 4394 20102 4406 20154
rect 4458 20102 4470 20154
rect 4522 20102 34934 20154
rect 34986 20102 34998 20154
rect 35050 20102 35062 20154
rect 35114 20102 35126 20154
rect 35178 20102 35190 20154
rect 35242 20102 58880 20154
rect 1104 20080 58880 20102
rect 1104 19610 58880 19632
rect 1104 19558 19574 19610
rect 19626 19558 19638 19610
rect 19690 19558 19702 19610
rect 19754 19558 19766 19610
rect 19818 19558 19830 19610
rect 19882 19558 50294 19610
rect 50346 19558 50358 19610
rect 50410 19558 50422 19610
rect 50474 19558 50486 19610
rect 50538 19558 50550 19610
rect 50602 19558 58880 19610
rect 1104 19536 58880 19558
rect 56134 19320 56140 19372
rect 56192 19360 56198 19372
rect 56321 19363 56379 19369
rect 56321 19360 56333 19363
rect 56192 19332 56333 19360
rect 56192 19320 56198 19332
rect 56321 19329 56333 19332
rect 56367 19329 56379 19363
rect 56321 19323 56379 19329
rect 56413 19159 56471 19165
rect 56413 19125 56425 19159
rect 56459 19156 56471 19159
rect 56502 19156 56508 19168
rect 56459 19128 56508 19156
rect 56459 19125 56471 19128
rect 56413 19119 56471 19125
rect 56502 19116 56508 19128
rect 56560 19116 56566 19168
rect 57882 19156 57888 19168
rect 57843 19128 57888 19156
rect 57882 19116 57888 19128
rect 57940 19116 57946 19168
rect 1104 19066 58880 19088
rect 1104 19014 4214 19066
rect 4266 19014 4278 19066
rect 4330 19014 4342 19066
rect 4394 19014 4406 19066
rect 4458 19014 4470 19066
rect 4522 19014 34934 19066
rect 34986 19014 34998 19066
rect 35050 19014 35062 19066
rect 35114 19014 35126 19066
rect 35178 19014 35190 19066
rect 35242 19014 58880 19066
rect 1104 18992 58880 19014
rect 57882 18884 57888 18896
rect 56336 18856 57888 18884
rect 56336 18825 56364 18856
rect 57882 18844 57888 18856
rect 57940 18844 57946 18896
rect 56321 18819 56379 18825
rect 56321 18785 56333 18819
rect 56367 18785 56379 18819
rect 56502 18816 56508 18828
rect 56463 18788 56508 18816
rect 56321 18779 56379 18785
rect 56502 18776 56508 18788
rect 56560 18776 56566 18828
rect 58158 18816 58164 18828
rect 58119 18788 58164 18816
rect 58158 18776 58164 18788
rect 58216 18776 58222 18828
rect 1104 18522 58880 18544
rect 1104 18470 19574 18522
rect 19626 18470 19638 18522
rect 19690 18470 19702 18522
rect 19754 18470 19766 18522
rect 19818 18470 19830 18522
rect 19882 18470 50294 18522
rect 50346 18470 50358 18522
rect 50410 18470 50422 18522
rect 50474 18470 50486 18522
rect 50538 18470 50550 18522
rect 50602 18470 58880 18522
rect 1104 18448 58880 18470
rect 1104 17978 58880 18000
rect 1104 17926 4214 17978
rect 4266 17926 4278 17978
rect 4330 17926 4342 17978
rect 4394 17926 4406 17978
rect 4458 17926 4470 17978
rect 4522 17926 34934 17978
rect 34986 17926 34998 17978
rect 35050 17926 35062 17978
rect 35114 17926 35126 17978
rect 35178 17926 35190 17978
rect 35242 17926 58880 17978
rect 1104 17904 58880 17926
rect 1104 17434 58880 17456
rect 1104 17382 19574 17434
rect 19626 17382 19638 17434
rect 19690 17382 19702 17434
rect 19754 17382 19766 17434
rect 19818 17382 19830 17434
rect 19882 17382 50294 17434
rect 50346 17382 50358 17434
rect 50410 17382 50422 17434
rect 50474 17382 50486 17434
rect 50538 17382 50550 17434
rect 50602 17382 58880 17434
rect 1104 17360 58880 17382
rect 1104 16890 58880 16912
rect 1104 16838 4214 16890
rect 4266 16838 4278 16890
rect 4330 16838 4342 16890
rect 4394 16838 4406 16890
rect 4458 16838 4470 16890
rect 4522 16838 34934 16890
rect 34986 16838 34998 16890
rect 35050 16838 35062 16890
rect 35114 16838 35126 16890
rect 35178 16838 35190 16890
rect 35242 16838 58880 16890
rect 1104 16816 58880 16838
rect 1104 16346 58880 16368
rect 1104 16294 19574 16346
rect 19626 16294 19638 16346
rect 19690 16294 19702 16346
rect 19754 16294 19766 16346
rect 19818 16294 19830 16346
rect 19882 16294 50294 16346
rect 50346 16294 50358 16346
rect 50410 16294 50422 16346
rect 50474 16294 50486 16346
rect 50538 16294 50550 16346
rect 50602 16294 58880 16346
rect 1104 16272 58880 16294
rect 1104 15802 58880 15824
rect 1104 15750 4214 15802
rect 4266 15750 4278 15802
rect 4330 15750 4342 15802
rect 4394 15750 4406 15802
rect 4458 15750 4470 15802
rect 4522 15750 34934 15802
rect 34986 15750 34998 15802
rect 35050 15750 35062 15802
rect 35114 15750 35126 15802
rect 35178 15750 35190 15802
rect 35242 15750 58880 15802
rect 1104 15728 58880 15750
rect 1104 15258 58880 15280
rect 1104 15206 19574 15258
rect 19626 15206 19638 15258
rect 19690 15206 19702 15258
rect 19754 15206 19766 15258
rect 19818 15206 19830 15258
rect 19882 15206 50294 15258
rect 50346 15206 50358 15258
rect 50410 15206 50422 15258
rect 50474 15206 50486 15258
rect 50538 15206 50550 15258
rect 50602 15206 58880 15258
rect 1104 15184 58880 15206
rect 1104 14714 58880 14736
rect 1104 14662 4214 14714
rect 4266 14662 4278 14714
rect 4330 14662 4342 14714
rect 4394 14662 4406 14714
rect 4458 14662 4470 14714
rect 4522 14662 34934 14714
rect 34986 14662 34998 14714
rect 35050 14662 35062 14714
rect 35114 14662 35126 14714
rect 35178 14662 35190 14714
rect 35242 14662 58880 14714
rect 1104 14640 58880 14662
rect 1104 14170 58880 14192
rect 1104 14118 19574 14170
rect 19626 14118 19638 14170
rect 19690 14118 19702 14170
rect 19754 14118 19766 14170
rect 19818 14118 19830 14170
rect 19882 14118 50294 14170
rect 50346 14118 50358 14170
rect 50410 14118 50422 14170
rect 50474 14118 50486 14170
rect 50538 14118 50550 14170
rect 50602 14118 58880 14170
rect 1104 14096 58880 14118
rect 1104 13626 58880 13648
rect 1104 13574 4214 13626
rect 4266 13574 4278 13626
rect 4330 13574 4342 13626
rect 4394 13574 4406 13626
rect 4458 13574 4470 13626
rect 4522 13574 34934 13626
rect 34986 13574 34998 13626
rect 35050 13574 35062 13626
rect 35114 13574 35126 13626
rect 35178 13574 35190 13626
rect 35242 13574 58880 13626
rect 1104 13552 58880 13574
rect 1104 13082 58880 13104
rect 1104 13030 19574 13082
rect 19626 13030 19638 13082
rect 19690 13030 19702 13082
rect 19754 13030 19766 13082
rect 19818 13030 19830 13082
rect 19882 13030 50294 13082
rect 50346 13030 50358 13082
rect 50410 13030 50422 13082
rect 50474 13030 50486 13082
rect 50538 13030 50550 13082
rect 50602 13030 58880 13082
rect 1104 13008 58880 13030
rect 1104 12538 58880 12560
rect 1104 12486 4214 12538
rect 4266 12486 4278 12538
rect 4330 12486 4342 12538
rect 4394 12486 4406 12538
rect 4458 12486 4470 12538
rect 4522 12486 34934 12538
rect 34986 12486 34998 12538
rect 35050 12486 35062 12538
rect 35114 12486 35126 12538
rect 35178 12486 35190 12538
rect 35242 12486 58880 12538
rect 1104 12464 58880 12486
rect 56318 12180 56324 12232
rect 56376 12220 56382 12232
rect 57241 12223 57299 12229
rect 57241 12220 57253 12223
rect 56376 12192 57253 12220
rect 56376 12180 56382 12192
rect 57241 12189 57253 12192
rect 57287 12189 57299 12223
rect 57241 12183 57299 12189
rect 1104 11994 58880 12016
rect 1104 11942 19574 11994
rect 19626 11942 19638 11994
rect 19690 11942 19702 11994
rect 19754 11942 19766 11994
rect 19818 11942 19830 11994
rect 19882 11942 50294 11994
rect 50346 11942 50358 11994
rect 50410 11942 50422 11994
rect 50474 11942 50486 11994
rect 50538 11942 50550 11994
rect 50602 11942 58880 11994
rect 1104 11920 58880 11942
rect 56962 11744 56968 11756
rect 56923 11716 56968 11744
rect 56962 11704 56968 11716
rect 57020 11704 57026 11756
rect 56502 11500 56508 11552
rect 56560 11540 56566 11552
rect 57057 11543 57115 11549
rect 57057 11540 57069 11543
rect 56560 11512 57069 11540
rect 56560 11500 56566 11512
rect 57057 11509 57069 11512
rect 57103 11509 57115 11543
rect 57057 11503 57115 11509
rect 1104 11450 58880 11472
rect 1104 11398 4214 11450
rect 4266 11398 4278 11450
rect 4330 11398 4342 11450
rect 4394 11398 4406 11450
rect 4458 11398 4470 11450
rect 4522 11398 34934 11450
rect 34986 11398 34998 11450
rect 35050 11398 35062 11450
rect 35114 11398 35126 11450
rect 35178 11398 35190 11450
rect 35242 11398 58880 11450
rect 1104 11376 58880 11398
rect 56318 11200 56324 11212
rect 56279 11172 56324 11200
rect 56318 11160 56324 11172
rect 56376 11160 56382 11212
rect 56502 11200 56508 11212
rect 56463 11172 56508 11200
rect 56502 11160 56508 11172
rect 56560 11160 56566 11212
rect 58158 11200 58164 11212
rect 58119 11172 58164 11200
rect 58158 11160 58164 11172
rect 58216 11160 58222 11212
rect 2501 11135 2559 11141
rect 2501 11101 2513 11135
rect 2547 11132 2559 11135
rect 8846 11132 8852 11144
rect 2547 11104 8852 11132
rect 2547 11101 2559 11104
rect 2501 11095 2559 11101
rect 8846 11092 8852 11104
rect 8904 11092 8910 11144
rect 2130 10956 2136 11008
rect 2188 10996 2194 11008
rect 2409 10999 2467 11005
rect 2409 10996 2421 10999
rect 2188 10968 2421 10996
rect 2188 10956 2194 10968
rect 2409 10965 2421 10968
rect 2455 10965 2467 10999
rect 2409 10959 2467 10965
rect 1104 10906 58880 10928
rect 1104 10854 19574 10906
rect 19626 10854 19638 10906
rect 19690 10854 19702 10906
rect 19754 10854 19766 10906
rect 19818 10854 19830 10906
rect 19882 10854 50294 10906
rect 50346 10854 50358 10906
rect 50410 10854 50422 10906
rect 50474 10854 50486 10906
rect 50538 10854 50550 10906
rect 50602 10854 58880 10906
rect 1104 10832 58880 10854
rect 2130 10724 2136 10736
rect 2091 10696 2136 10724
rect 2130 10684 2136 10696
rect 2188 10684 2194 10736
rect 1946 10588 1952 10600
rect 1907 10560 1952 10588
rect 1946 10548 1952 10560
rect 2004 10548 2010 10600
rect 2774 10588 2780 10600
rect 2735 10560 2780 10588
rect 2774 10548 2780 10560
rect 2832 10548 2838 10600
rect 1104 10362 58880 10384
rect 1104 10310 4214 10362
rect 4266 10310 4278 10362
rect 4330 10310 4342 10362
rect 4394 10310 4406 10362
rect 4458 10310 4470 10362
rect 4522 10310 34934 10362
rect 34986 10310 34998 10362
rect 35050 10310 35062 10362
rect 35114 10310 35126 10362
rect 35178 10310 35190 10362
rect 35242 10310 58880 10362
rect 1104 10288 58880 10310
rect 1946 10208 1952 10260
rect 2004 10248 2010 10260
rect 2041 10251 2099 10257
rect 2041 10248 2053 10251
rect 2004 10220 2053 10248
rect 2004 10208 2010 10220
rect 2041 10217 2053 10220
rect 2087 10217 2099 10251
rect 2041 10211 2099 10217
rect 1104 9818 58880 9840
rect 1104 9766 19574 9818
rect 19626 9766 19638 9818
rect 19690 9766 19702 9818
rect 19754 9766 19766 9818
rect 19818 9766 19830 9818
rect 19882 9766 50294 9818
rect 50346 9766 50358 9818
rect 50410 9766 50422 9818
rect 50474 9766 50486 9818
rect 50538 9766 50550 9818
rect 50602 9766 58880 9818
rect 1104 9744 58880 9766
rect 1104 9274 58880 9296
rect 1104 9222 4214 9274
rect 4266 9222 4278 9274
rect 4330 9222 4342 9274
rect 4394 9222 4406 9274
rect 4458 9222 4470 9274
rect 4522 9222 34934 9274
rect 34986 9222 34998 9274
rect 35050 9222 35062 9274
rect 35114 9222 35126 9274
rect 35178 9222 35190 9274
rect 35242 9222 58880 9274
rect 1104 9200 58880 9222
rect 56321 9027 56379 9033
rect 56321 8993 56333 9027
rect 56367 9024 56379 9027
rect 57882 9024 57888 9036
rect 56367 8996 57888 9024
rect 56367 8993 56379 8996
rect 56321 8987 56379 8993
rect 57882 8984 57888 8996
rect 57940 8984 57946 9036
rect 56502 8888 56508 8900
rect 56463 8860 56508 8888
rect 56502 8848 56508 8860
rect 56560 8848 56566 8900
rect 58158 8888 58164 8900
rect 58119 8860 58164 8888
rect 58158 8848 58164 8860
rect 58216 8848 58222 8900
rect 1104 8730 58880 8752
rect 1104 8678 19574 8730
rect 19626 8678 19638 8730
rect 19690 8678 19702 8730
rect 19754 8678 19766 8730
rect 19818 8678 19830 8730
rect 19882 8678 50294 8730
rect 50346 8678 50358 8730
rect 50410 8678 50422 8730
rect 50474 8678 50486 8730
rect 50538 8678 50550 8730
rect 50602 8678 58880 8730
rect 1104 8656 58880 8678
rect 56413 8619 56471 8625
rect 56413 8585 56425 8619
rect 56459 8616 56471 8619
rect 56502 8616 56508 8628
rect 56459 8588 56508 8616
rect 56459 8585 56471 8588
rect 56413 8579 56471 8585
rect 56502 8576 56508 8588
rect 56560 8576 56566 8628
rect 56226 8440 56232 8492
rect 56284 8480 56290 8492
rect 56321 8483 56379 8489
rect 56321 8480 56333 8483
rect 56284 8452 56333 8480
rect 56284 8440 56290 8452
rect 56321 8449 56333 8452
rect 56367 8449 56379 8483
rect 57882 8480 57888 8492
rect 57843 8452 57888 8480
rect 56321 8443 56379 8449
rect 57882 8440 57888 8452
rect 57940 8440 57946 8492
rect 1104 8186 58880 8208
rect 1104 8134 4214 8186
rect 4266 8134 4278 8186
rect 4330 8134 4342 8186
rect 4394 8134 4406 8186
rect 4458 8134 4470 8186
rect 4522 8134 34934 8186
rect 34986 8134 34998 8186
rect 35050 8134 35062 8186
rect 35114 8134 35126 8186
rect 35178 8134 35190 8186
rect 35242 8134 58880 8186
rect 1104 8112 58880 8134
rect 1104 7642 58880 7664
rect 1104 7590 19574 7642
rect 19626 7590 19638 7642
rect 19690 7590 19702 7642
rect 19754 7590 19766 7642
rect 19818 7590 19830 7642
rect 19882 7590 50294 7642
rect 50346 7590 50358 7642
rect 50410 7590 50422 7642
rect 50474 7590 50486 7642
rect 50538 7590 50550 7642
rect 50602 7590 58880 7642
rect 1104 7568 58880 7590
rect 1104 7098 58880 7120
rect 1104 7046 4214 7098
rect 4266 7046 4278 7098
rect 4330 7046 4342 7098
rect 4394 7046 4406 7098
rect 4458 7046 4470 7098
rect 4522 7046 34934 7098
rect 34986 7046 34998 7098
rect 35050 7046 35062 7098
rect 35114 7046 35126 7098
rect 35178 7046 35190 7098
rect 35242 7046 58880 7098
rect 1104 7024 58880 7046
rect 1104 6554 58880 6576
rect 1104 6502 19574 6554
rect 19626 6502 19638 6554
rect 19690 6502 19702 6554
rect 19754 6502 19766 6554
rect 19818 6502 19830 6554
rect 19882 6502 50294 6554
rect 50346 6502 50358 6554
rect 50410 6502 50422 6554
rect 50474 6502 50486 6554
rect 50538 6502 50550 6554
rect 50602 6502 58880 6554
rect 1104 6480 58880 6502
rect 1104 6010 58880 6032
rect 1104 5958 4214 6010
rect 4266 5958 4278 6010
rect 4330 5958 4342 6010
rect 4394 5958 4406 6010
rect 4458 5958 4470 6010
rect 4522 5958 34934 6010
rect 34986 5958 34998 6010
rect 35050 5958 35062 6010
rect 35114 5958 35126 6010
rect 35178 5958 35190 6010
rect 35242 5958 58880 6010
rect 1104 5936 58880 5958
rect 1104 5466 58880 5488
rect 1104 5414 19574 5466
rect 19626 5414 19638 5466
rect 19690 5414 19702 5466
rect 19754 5414 19766 5466
rect 19818 5414 19830 5466
rect 19882 5414 50294 5466
rect 50346 5414 50358 5466
rect 50410 5414 50422 5466
rect 50474 5414 50486 5466
rect 50538 5414 50550 5466
rect 50602 5414 58880 5466
rect 1104 5392 58880 5414
rect 1946 4972 1952 5024
rect 2004 5012 2010 5024
rect 2041 5015 2099 5021
rect 2041 5012 2053 5015
rect 2004 4984 2053 5012
rect 2004 4972 2010 4984
rect 2041 4981 2053 4984
rect 2087 4981 2099 5015
rect 2041 4975 2099 4981
rect 1104 4922 58880 4944
rect 1104 4870 4214 4922
rect 4266 4870 4278 4922
rect 4330 4870 4342 4922
rect 4394 4870 4406 4922
rect 4458 4870 4470 4922
rect 4522 4870 34934 4922
rect 34986 4870 34998 4922
rect 35050 4870 35062 4922
rect 35114 4870 35126 4922
rect 35178 4870 35190 4922
rect 35242 4870 58880 4922
rect 1104 4848 58880 4870
rect 2498 4604 2504 4616
rect 2411 4576 2504 4604
rect 2498 4564 2504 4576
rect 2556 4604 2562 4616
rect 8202 4604 8208 4616
rect 2556 4576 8208 4604
rect 2556 4564 2562 4576
rect 8202 4564 8208 4576
rect 8260 4564 8266 4616
rect 56318 4604 56324 4616
rect 56279 4576 56324 4604
rect 56318 4564 56324 4576
rect 56376 4564 56382 4616
rect 56502 4536 56508 4548
rect 56463 4508 56508 4536
rect 56502 4496 56508 4508
rect 56560 4496 56566 4548
rect 58161 4539 58219 4545
rect 58161 4505 58173 4539
rect 58207 4536 58219 4539
rect 59262 4536 59268 4548
rect 58207 4508 59268 4536
rect 58207 4505 58219 4508
rect 58161 4499 58219 4505
rect 59262 4496 59268 4508
rect 59320 4496 59326 4548
rect 2130 4428 2136 4480
rect 2188 4468 2194 4480
rect 2409 4471 2467 4477
rect 2409 4468 2421 4471
rect 2188 4440 2421 4468
rect 2188 4428 2194 4440
rect 2409 4437 2421 4440
rect 2455 4437 2467 4471
rect 2409 4431 2467 4437
rect 1104 4378 58880 4400
rect 1104 4326 19574 4378
rect 19626 4326 19638 4378
rect 19690 4326 19702 4378
rect 19754 4326 19766 4378
rect 19818 4326 19830 4378
rect 19882 4326 50294 4378
rect 50346 4326 50358 4378
rect 50410 4326 50422 4378
rect 50474 4326 50486 4378
rect 50538 4326 50550 4378
rect 50602 4326 58880 4378
rect 1104 4304 58880 4326
rect 2130 4196 2136 4208
rect 2091 4168 2136 4196
rect 2130 4156 2136 4168
rect 2188 4156 2194 4208
rect 1946 4128 1952 4140
rect 1907 4100 1952 4128
rect 1946 4088 1952 4100
rect 2004 4088 2010 4140
rect 7558 4128 7564 4140
rect 7519 4100 7564 4128
rect 7558 4088 7564 4100
rect 7616 4088 7622 4140
rect 57790 4088 57796 4140
rect 57848 4128 57854 4140
rect 57885 4131 57943 4137
rect 57885 4128 57897 4131
rect 57848 4100 57897 4128
rect 57848 4088 57854 4100
rect 57885 4097 57897 4100
rect 57931 4097 57943 4131
rect 57885 4091 57943 4097
rect 2774 4060 2780 4072
rect 2735 4032 2780 4060
rect 2774 4020 2780 4032
rect 2832 4020 2838 4072
rect 4706 4020 4712 4072
rect 4764 4060 4770 4072
rect 8757 4063 8815 4069
rect 8757 4060 8769 4063
rect 4764 4032 8769 4060
rect 4764 4020 4770 4032
rect 8757 4029 8769 4032
rect 8803 4060 8815 4063
rect 51442 4060 51448 4072
rect 8803 4032 51448 4060
rect 8803 4029 8815 4032
rect 8757 4023 8815 4029
rect 51442 4020 51448 4032
rect 51500 4020 51506 4072
rect 56873 4063 56931 4069
rect 56873 4029 56885 4063
rect 56919 4029 56931 4063
rect 56873 4023 56931 4029
rect 57149 4063 57207 4069
rect 57149 4029 57161 4063
rect 57195 4029 57207 4063
rect 57330 4060 57336 4072
rect 57291 4032 57336 4060
rect 57149 4023 57207 4029
rect 4062 3884 4068 3936
rect 4120 3924 4126 3936
rect 4249 3927 4307 3933
rect 4249 3924 4261 3927
rect 4120 3896 4261 3924
rect 4120 3884 4126 3896
rect 4249 3893 4261 3896
rect 4295 3893 4307 3927
rect 4249 3887 4307 3893
rect 20622 3884 20628 3936
rect 20680 3924 20686 3936
rect 20717 3927 20775 3933
rect 20717 3924 20729 3927
rect 20680 3896 20729 3924
rect 20680 3884 20686 3896
rect 20717 3893 20729 3896
rect 20763 3893 20775 3927
rect 51534 3924 51540 3936
rect 51495 3896 51540 3924
rect 20717 3887 20775 3893
rect 51534 3884 51540 3896
rect 51592 3884 51598 3936
rect 54478 3924 54484 3936
rect 54439 3896 54484 3924
rect 54478 3884 54484 3896
rect 54536 3884 54542 3936
rect 56888 3924 56916 4023
rect 57164 3992 57192 4023
rect 57330 4020 57336 4032
rect 57388 4020 57394 4072
rect 57977 3995 58035 4001
rect 57977 3992 57989 3995
rect 57164 3964 57989 3992
rect 57977 3961 57989 3964
rect 58023 3961 58035 3995
rect 57977 3955 58035 3961
rect 57238 3924 57244 3936
rect 56888 3896 57244 3924
rect 57238 3884 57244 3896
rect 57296 3884 57302 3936
rect 1104 3834 58880 3856
rect 1104 3782 4214 3834
rect 4266 3782 4278 3834
rect 4330 3782 4342 3834
rect 4394 3782 4406 3834
rect 4458 3782 4470 3834
rect 4522 3782 34934 3834
rect 34986 3782 34998 3834
rect 35050 3782 35062 3834
rect 35114 3782 35126 3834
rect 35178 3782 35190 3834
rect 35242 3782 58880 3834
rect 1104 3760 58880 3782
rect 55769 3723 55827 3729
rect 55769 3689 55781 3723
rect 55815 3720 55827 3723
rect 56502 3720 56508 3732
rect 55815 3692 56508 3720
rect 55815 3689 55827 3692
rect 55769 3683 55827 3689
rect 56502 3680 56508 3692
rect 56560 3680 56566 3732
rect 56778 3652 56784 3664
rect 44284 3624 56784 3652
rect 4062 3584 4068 3596
rect 4023 3556 4068 3584
rect 4062 3544 4068 3556
rect 4120 3544 4126 3596
rect 4614 3584 4620 3596
rect 4575 3556 4620 3584
rect 4614 3544 4620 3556
rect 4672 3544 4678 3596
rect 14182 3544 14188 3596
rect 14240 3584 14246 3596
rect 14921 3587 14979 3593
rect 14921 3584 14933 3587
rect 14240 3556 14933 3584
rect 14240 3544 14246 3556
rect 14921 3553 14933 3556
rect 14967 3553 14979 3587
rect 14921 3547 14979 3553
rect 16546 3556 26234 3584
rect 7558 3516 7564 3528
rect 7519 3488 7564 3516
rect 7558 3476 7564 3488
rect 7616 3476 7622 3528
rect 14458 3516 14464 3528
rect 14419 3488 14464 3516
rect 14458 3476 14464 3488
rect 14516 3476 14522 3528
rect 4246 3448 4252 3460
rect 4207 3420 4252 3448
rect 4246 3408 4252 3420
rect 4304 3408 4310 3460
rect 8202 3448 8208 3460
rect 8115 3420 8208 3448
rect 8202 3408 8208 3420
rect 8260 3408 8266 3460
rect 14645 3451 14703 3457
rect 14645 3417 14657 3451
rect 14691 3448 14703 3451
rect 15470 3448 15476 3460
rect 14691 3420 15476 3448
rect 14691 3417 14703 3420
rect 14645 3411 14703 3417
rect 15470 3408 15476 3420
rect 15528 3408 15534 3460
rect 8220 3380 8248 3408
rect 16546 3380 16574 3556
rect 18690 3476 18696 3528
rect 18748 3516 18754 3528
rect 20622 3516 20628 3528
rect 18748 3488 18793 3516
rect 20583 3488 20628 3516
rect 18748 3476 18754 3488
rect 20622 3476 20628 3488
rect 20680 3476 20686 3528
rect 26206 3516 26234 3556
rect 44284 3525 44312 3624
rect 56778 3612 56784 3624
rect 56836 3612 56842 3664
rect 45186 3544 45192 3596
rect 45244 3584 45250 3596
rect 45465 3587 45523 3593
rect 45465 3584 45477 3587
rect 45244 3556 45477 3584
rect 45244 3544 45250 3556
rect 45465 3553 45477 3556
rect 45511 3553 45523 3587
rect 51534 3584 51540 3596
rect 51495 3556 51540 3584
rect 45465 3547 45523 3553
rect 51534 3544 51540 3556
rect 51592 3544 51598 3596
rect 52178 3584 52184 3596
rect 52139 3556 52184 3584
rect 52178 3544 52184 3556
rect 52236 3544 52242 3596
rect 57882 3584 57888 3596
rect 57843 3556 57888 3584
rect 57882 3544 57888 3556
rect 57940 3544 57946 3596
rect 44269 3519 44327 3525
rect 44269 3516 44281 3519
rect 26206 3488 44281 3516
rect 44269 3485 44281 3488
rect 44315 3485 44327 3519
rect 44269 3479 44327 3485
rect 44634 3476 44640 3528
rect 44692 3516 44698 3528
rect 45005 3519 45063 3525
rect 45005 3516 45017 3519
rect 44692 3488 45017 3516
rect 44692 3476 44698 3488
rect 45005 3485 45017 3488
rect 45051 3485 45063 3519
rect 54573 3519 54631 3525
rect 54573 3516 54585 3519
rect 45005 3479 45063 3485
rect 52932 3488 54585 3516
rect 16758 3408 16764 3460
rect 16816 3448 16822 3460
rect 16853 3451 16911 3457
rect 16853 3448 16865 3451
rect 16816 3420 16865 3448
rect 16816 3408 16822 3420
rect 16853 3417 16865 3420
rect 16899 3417 16911 3451
rect 16853 3411 16911 3417
rect 18414 3408 18420 3460
rect 18472 3448 18478 3460
rect 18509 3451 18567 3457
rect 18509 3448 18521 3451
rect 18472 3420 18521 3448
rect 18472 3408 18478 3420
rect 18509 3417 18521 3420
rect 18555 3417 18567 3451
rect 20806 3448 20812 3460
rect 20767 3420 20812 3448
rect 18509 3411 18567 3417
rect 20806 3408 20812 3420
rect 20864 3408 20870 3460
rect 21266 3408 21272 3460
rect 21324 3448 21330 3460
rect 22465 3451 22523 3457
rect 22465 3448 22477 3451
rect 21324 3420 22477 3448
rect 21324 3408 21330 3420
rect 22465 3417 22477 3420
rect 22511 3417 22523 3451
rect 22465 3411 22523 3417
rect 44361 3451 44419 3457
rect 44361 3417 44373 3451
rect 44407 3448 44419 3451
rect 45189 3451 45247 3457
rect 45189 3448 45201 3451
rect 44407 3420 45201 3448
rect 44407 3417 44419 3420
rect 44361 3411 44419 3417
rect 45189 3417 45201 3420
rect 45235 3417 45247 3451
rect 51718 3448 51724 3460
rect 51679 3420 51724 3448
rect 45189 3411 45247 3417
rect 51718 3408 51724 3420
rect 51776 3408 51782 3460
rect 8220 3352 16574 3380
rect 50154 3340 50160 3392
rect 50212 3380 50218 3392
rect 52932 3380 52960 3488
rect 54573 3485 54585 3488
rect 54619 3516 54631 3519
rect 55674 3516 55680 3528
rect 54619 3488 55680 3516
rect 54619 3485 54631 3488
rect 54573 3479 54631 3485
rect 55674 3476 55680 3488
rect 55732 3476 55738 3528
rect 56318 3516 56324 3528
rect 56279 3488 56324 3516
rect 56318 3476 56324 3488
rect 56376 3476 56382 3528
rect 56505 3451 56563 3457
rect 56505 3417 56517 3451
rect 56551 3448 56563 3451
rect 56870 3448 56876 3460
rect 56551 3420 56876 3448
rect 56551 3417 56563 3420
rect 56505 3411 56563 3417
rect 56870 3408 56876 3420
rect 56928 3408 56934 3460
rect 54662 3380 54668 3392
rect 50212 3352 52960 3380
rect 54623 3352 54668 3380
rect 50212 3340 50218 3352
rect 54662 3340 54668 3352
rect 54720 3340 54726 3392
rect 1104 3290 58880 3312
rect 1104 3238 19574 3290
rect 19626 3238 19638 3290
rect 19690 3238 19702 3290
rect 19754 3238 19766 3290
rect 19818 3238 19830 3290
rect 19882 3238 50294 3290
rect 50346 3238 50358 3290
rect 50410 3238 50422 3290
rect 50474 3238 50486 3290
rect 50538 3238 50550 3290
rect 50602 3238 58880 3290
rect 1104 3216 58880 3238
rect 4246 3176 4252 3188
rect 4207 3148 4252 3176
rect 4246 3136 4252 3148
rect 4304 3136 4310 3188
rect 15470 3176 15476 3188
rect 15431 3148 15476 3176
rect 15470 3136 15476 3148
rect 15528 3136 15534 3188
rect 18414 3176 18420 3188
rect 18375 3148 18420 3176
rect 18414 3136 18420 3148
rect 18472 3136 18478 3188
rect 20806 3176 20812 3188
rect 20767 3148 20812 3176
rect 20806 3136 20812 3148
rect 20864 3136 20870 3188
rect 51629 3179 51687 3185
rect 51629 3145 51641 3179
rect 51675 3176 51687 3179
rect 51718 3176 51724 3188
rect 51675 3148 51724 3176
rect 51675 3145 51687 3148
rect 51629 3139 51687 3145
rect 51718 3136 51724 3148
rect 51776 3136 51782 3188
rect 56134 3176 56140 3188
rect 51828 3148 56140 3176
rect 18690 3108 18696 3120
rect 17420 3080 18696 3108
rect 4157 3043 4215 3049
rect 4157 3009 4169 3043
rect 4203 3040 4215 3043
rect 4706 3040 4712 3052
rect 4203 3012 4712 3040
rect 4203 3009 4215 3012
rect 4157 3003 4215 3009
rect 4706 3000 4712 3012
rect 4764 3000 4770 3052
rect 14458 3040 14464 3052
rect 14419 3012 14464 3040
rect 14458 3000 14464 3012
rect 14516 3000 14522 3052
rect 17420 3049 17448 3080
rect 18690 3068 18696 3080
rect 18748 3068 18754 3120
rect 51828 3108 51856 3148
rect 56134 3136 56140 3148
rect 56192 3136 56198 3188
rect 56870 3176 56876 3188
rect 56831 3148 56876 3176
rect 56870 3136 56876 3148
rect 56928 3136 56934 3188
rect 54662 3108 54668 3120
rect 26206 3080 50384 3108
rect 15565 3043 15623 3049
rect 15565 3009 15577 3043
rect 15611 3040 15623 3043
rect 17405 3043 17463 3049
rect 15611 3012 16574 3040
rect 15611 3009 15623 3012
rect 15565 3003 15623 3009
rect 16546 2904 16574 3012
rect 17405 3009 17417 3043
rect 17451 3009 17463 3043
rect 17405 3003 17463 3009
rect 18509 3043 18567 3049
rect 18509 3009 18521 3043
rect 18555 3040 18567 3043
rect 20717 3043 20775 3049
rect 20717 3040 20729 3043
rect 18555 3012 20729 3040
rect 18555 3009 18567 3012
rect 18509 3003 18567 3009
rect 20717 3009 20729 3012
rect 20763 3040 20775 3043
rect 26206 3040 26234 3080
rect 44634 3040 44640 3052
rect 20763 3012 26234 3040
rect 44595 3012 44640 3040
rect 20763 3009 20775 3012
rect 20717 3003 20775 3009
rect 44634 3000 44640 3012
rect 44692 3000 44698 3052
rect 50154 2904 50160 2916
rect 16546 2876 50160 2904
rect 50154 2864 50160 2876
rect 50212 2864 50218 2916
rect 50356 2904 50384 3080
rect 51552 3080 51856 3108
rect 54623 3080 54668 3108
rect 51442 3000 51448 3052
rect 51500 3040 51506 3052
rect 51552 3049 51580 3080
rect 54662 3068 54668 3080
rect 54720 3068 54726 3120
rect 56318 3068 56324 3120
rect 56376 3108 56382 3120
rect 56376 3080 57928 3108
rect 56376 3068 56382 3080
rect 51537 3043 51595 3049
rect 51537 3040 51549 3043
rect 51500 3012 51549 3040
rect 51500 3000 51506 3012
rect 51537 3009 51549 3012
rect 51583 3009 51595 3043
rect 54478 3040 54484 3052
rect 54439 3012 54484 3040
rect 51537 3003 51595 3009
rect 54478 3000 54484 3012
rect 54536 3000 54542 3052
rect 56778 3040 56784 3052
rect 56739 3012 56784 3040
rect 56778 3000 56784 3012
rect 56836 3000 56842 3052
rect 57900 3049 57928 3080
rect 57885 3043 57943 3049
rect 57885 3009 57897 3043
rect 57931 3009 57943 3043
rect 57885 3003 57943 3009
rect 54754 2932 54760 2984
rect 54812 2972 54818 2984
rect 54941 2975 54999 2981
rect 54941 2972 54953 2975
rect 54812 2944 54953 2972
rect 54812 2932 54818 2944
rect 54941 2941 54953 2944
rect 54987 2941 54999 2975
rect 54941 2935 54999 2941
rect 56226 2904 56232 2916
rect 50356 2876 56232 2904
rect 56226 2864 56232 2876
rect 56284 2864 56290 2916
rect 1104 2746 58880 2768
rect 1104 2694 4214 2746
rect 4266 2694 4278 2746
rect 4330 2694 4342 2746
rect 4394 2694 4406 2746
rect 4458 2694 4470 2746
rect 4522 2694 34934 2746
rect 34986 2694 34998 2746
rect 35050 2694 35062 2746
rect 35114 2694 35126 2746
rect 35178 2694 35190 2746
rect 35242 2694 58880 2746
rect 1104 2672 58880 2694
rect 7558 2632 7564 2644
rect 7519 2604 7564 2632
rect 7558 2592 7564 2604
rect 7616 2592 7622 2644
rect 56781 2635 56839 2641
rect 56781 2601 56793 2635
rect 56827 2632 56839 2635
rect 57330 2632 57336 2644
rect 56827 2604 57336 2632
rect 56827 2601 56839 2604
rect 56781 2595 56839 2601
rect 57330 2592 57336 2604
rect 57388 2592 57394 2644
rect 56410 2524 56416 2576
rect 56468 2564 56474 2576
rect 57885 2567 57943 2573
rect 57885 2564 57897 2567
rect 56468 2536 57897 2564
rect 56468 2524 56474 2536
rect 57885 2533 57897 2536
rect 57931 2533 57943 2567
rect 57885 2527 57943 2533
rect 23842 2388 23848 2440
rect 23900 2428 23906 2440
rect 24489 2431 24547 2437
rect 24489 2428 24501 2431
rect 23900 2400 24501 2428
rect 23900 2388 23906 2400
rect 24489 2397 24501 2400
rect 24535 2397 24547 2431
rect 24489 2391 24547 2397
rect 7098 2320 7104 2372
rect 7156 2360 7162 2372
rect 7285 2363 7343 2369
rect 7285 2360 7297 2363
rect 7156 2332 7297 2360
rect 7156 2320 7162 2332
rect 7285 2329 7297 2332
rect 7331 2329 7343 2363
rect 7285 2323 7343 2329
rect 25041 2363 25099 2369
rect 25041 2329 25053 2363
rect 25087 2360 25099 2363
rect 41506 2360 41512 2372
rect 25087 2332 41512 2360
rect 25087 2329 25099 2332
rect 25041 2323 25099 2329
rect 41506 2320 41512 2332
rect 41564 2320 41570 2372
rect 1104 2202 58880 2224
rect 1104 2150 19574 2202
rect 19626 2150 19638 2202
rect 19690 2150 19702 2202
rect 19754 2150 19766 2202
rect 19818 2150 19830 2202
rect 19882 2150 50294 2202
rect 50346 2150 50358 2202
rect 50410 2150 50422 2202
rect 50474 2150 50486 2202
rect 50538 2150 50550 2202
rect 50602 2150 58880 2202
rect 1104 2128 58880 2150
<< via1 >>
rect 19574 57638 19626 57690
rect 19638 57638 19690 57690
rect 19702 57638 19754 57690
rect 19766 57638 19818 57690
rect 19830 57638 19882 57690
rect 50294 57638 50346 57690
rect 50358 57638 50410 57690
rect 50422 57638 50474 57690
rect 50486 57638 50538 57690
rect 50550 57638 50602 57690
rect 41236 57400 41288 57452
rect 41696 57375 41748 57384
rect 41696 57341 41705 57375
rect 41705 57341 41739 57375
rect 41739 57341 41748 57375
rect 41696 57332 41748 57341
rect 4214 57094 4266 57146
rect 4278 57094 4330 57146
rect 4342 57094 4394 57146
rect 4406 57094 4458 57146
rect 4470 57094 4522 57146
rect 34934 57094 34986 57146
rect 34998 57094 35050 57146
rect 35062 57094 35114 57146
rect 35126 57094 35178 57146
rect 35190 57094 35242 57146
rect 8484 56788 8536 56840
rect 8944 56788 8996 56840
rect 25964 56788 26016 56840
rect 33508 56788 33560 56840
rect 35716 56831 35768 56840
rect 35716 56797 35725 56831
rect 35725 56797 35759 56831
rect 35759 56797 35768 56831
rect 35716 56788 35768 56797
rect 42524 56831 42576 56840
rect 42524 56797 42533 56831
rect 42533 56797 42567 56831
rect 42567 56797 42576 56831
rect 42524 56788 42576 56797
rect 43168 56831 43220 56840
rect 43168 56797 43177 56831
rect 43177 56797 43211 56831
rect 43211 56797 43220 56831
rect 43168 56788 43220 56797
rect 49884 56788 49936 56840
rect 52828 56788 52880 56840
rect 19574 56550 19626 56602
rect 19638 56550 19690 56602
rect 19702 56550 19754 56602
rect 19766 56550 19818 56602
rect 19830 56550 19882 56602
rect 50294 56550 50346 56602
rect 50358 56550 50410 56602
rect 50422 56550 50474 56602
rect 50486 56550 50538 56602
rect 50550 56550 50602 56602
rect 664 56380 716 56432
rect 8484 56355 8536 56364
rect 8484 56321 8493 56355
rect 8493 56321 8527 56355
rect 8527 56321 8536 56355
rect 8944 56355 8996 56364
rect 8484 56312 8536 56321
rect 8944 56321 8953 56355
rect 8953 56321 8987 56355
rect 8987 56321 8996 56355
rect 8944 56312 8996 56321
rect 33508 56355 33560 56364
rect 33508 56321 33517 56355
rect 33517 56321 33551 56355
rect 33551 56321 33560 56355
rect 33508 56312 33560 56321
rect 49884 56355 49936 56364
rect 49884 56321 49893 56355
rect 49893 56321 49927 56355
rect 49927 56321 49936 56355
rect 49884 56312 49936 56321
rect 52828 56355 52880 56364
rect 52828 56321 52837 56355
rect 52837 56321 52871 56355
rect 52871 56321 52880 56355
rect 52828 56312 52880 56321
rect 7748 56287 7800 56296
rect 7748 56253 7757 56287
rect 7757 56253 7791 56287
rect 7791 56253 7800 56287
rect 7748 56244 7800 56253
rect 8208 56244 8260 56296
rect 9128 56287 9180 56296
rect 9128 56253 9137 56287
rect 9137 56253 9171 56287
rect 9171 56253 9180 56287
rect 9128 56244 9180 56253
rect 9680 56287 9732 56296
rect 9680 56253 9689 56287
rect 9689 56253 9723 56287
rect 9723 56253 9732 56287
rect 9680 56244 9732 56253
rect 33692 56287 33744 56296
rect 33692 56253 33701 56287
rect 33701 56253 33735 56287
rect 33735 56253 33744 56287
rect 33692 56244 33744 56253
rect 34152 56287 34204 56296
rect 34152 56253 34161 56287
rect 34161 56253 34195 56287
rect 34195 56253 34204 56287
rect 34152 56244 34204 56253
rect 44364 56244 44416 56296
rect 45100 56287 45152 56296
rect 45100 56253 45109 56287
rect 45109 56253 45143 56287
rect 45143 56253 45152 56287
rect 45100 56244 45152 56253
rect 50252 56244 50304 56296
rect 50896 56244 50948 56296
rect 53196 56244 53248 56296
rect 26056 56176 26108 56228
rect 50344 56176 50396 56228
rect 52920 56176 52972 56228
rect 43720 56108 43772 56160
rect 4214 56006 4266 56058
rect 4278 56006 4330 56058
rect 4342 56006 4394 56058
rect 4406 56006 4458 56058
rect 4470 56006 4522 56058
rect 34934 56006 34986 56058
rect 34998 56006 35050 56058
rect 35062 56006 35114 56058
rect 35126 56006 35178 56058
rect 35190 56006 35242 56058
rect 33692 55947 33744 55956
rect 33692 55913 33701 55947
rect 33701 55913 33735 55947
rect 33735 55913 33744 55947
rect 33692 55904 33744 55913
rect 44364 55947 44416 55956
rect 25964 55811 26016 55820
rect 25964 55777 25973 55811
rect 25973 55777 26007 55811
rect 26007 55777 26016 55811
rect 25964 55768 26016 55777
rect 26424 55811 26476 55820
rect 26424 55777 26433 55811
rect 26433 55777 26467 55811
rect 26467 55777 26476 55811
rect 26424 55768 26476 55777
rect 35716 55811 35768 55820
rect 35716 55777 35725 55811
rect 35725 55777 35759 55811
rect 35759 55777 35768 55811
rect 35716 55768 35768 55777
rect 36084 55768 36136 55820
rect 41696 55768 41748 55820
rect 42524 55768 42576 55820
rect 44364 55913 44373 55947
rect 44373 55913 44407 55947
rect 44407 55913 44416 55947
rect 44364 55904 44416 55913
rect 50252 55947 50304 55956
rect 50252 55913 50261 55947
rect 50261 55913 50295 55947
rect 50295 55913 50304 55947
rect 50252 55904 50304 55913
rect 53196 55947 53248 55956
rect 53196 55913 53205 55947
rect 53205 55913 53239 55947
rect 53239 55913 53248 55947
rect 53196 55904 53248 55913
rect 33600 55743 33652 55752
rect 33600 55709 33609 55743
rect 33609 55709 33643 55743
rect 33643 55709 33652 55743
rect 33600 55700 33652 55709
rect 42708 55743 42760 55752
rect 42708 55709 42717 55743
rect 42717 55709 42751 55743
rect 42751 55709 42760 55743
rect 42708 55700 42760 55709
rect 43444 55700 43496 55752
rect 49700 55700 49752 55752
rect 50344 55745 50396 55752
rect 50344 55711 50361 55745
rect 50361 55711 50395 55745
rect 50395 55711 50396 55745
rect 50344 55700 50396 55711
rect 26148 55675 26200 55684
rect 26148 55641 26157 55675
rect 26157 55641 26191 55675
rect 26191 55641 26200 55675
rect 26148 55632 26200 55641
rect 35900 55675 35952 55684
rect 35900 55641 35909 55675
rect 35909 55641 35943 55675
rect 35943 55641 35952 55675
rect 56876 55700 56928 55752
rect 35900 55632 35952 55641
rect 55588 55632 55640 55684
rect 42984 55564 43036 55616
rect 43076 55564 43128 55616
rect 19574 55462 19626 55514
rect 19638 55462 19690 55514
rect 19702 55462 19754 55514
rect 19766 55462 19818 55514
rect 19830 55462 19882 55514
rect 50294 55462 50346 55514
rect 50358 55462 50410 55514
rect 50422 55462 50474 55514
rect 50486 55462 50538 55514
rect 50550 55462 50602 55514
rect 9128 55403 9180 55412
rect 9128 55369 9137 55403
rect 9137 55369 9171 55403
rect 9171 55369 9180 55403
rect 9128 55360 9180 55369
rect 26148 55403 26200 55412
rect 26148 55369 26157 55403
rect 26157 55369 26191 55403
rect 26191 55369 26200 55403
rect 26148 55360 26200 55369
rect 35900 55403 35952 55412
rect 35900 55369 35909 55403
rect 35909 55369 35943 55403
rect 35943 55369 35952 55403
rect 35900 55360 35952 55369
rect 42708 55360 42760 55412
rect 43536 55360 43588 55412
rect 49700 55360 49752 55412
rect 56232 55360 56284 55412
rect 9036 55267 9088 55276
rect 9036 55233 9045 55267
rect 9045 55233 9079 55267
rect 9079 55233 9088 55267
rect 9036 55224 9088 55233
rect 26056 55267 26108 55276
rect 26056 55233 26065 55267
rect 26065 55233 26099 55267
rect 26099 55233 26108 55267
rect 26056 55224 26108 55233
rect 43444 55224 43496 55276
rect 44180 55224 44232 55276
rect 43720 55156 43772 55208
rect 42340 55020 42392 55072
rect 4214 54918 4266 54970
rect 4278 54918 4330 54970
rect 4342 54918 4394 54970
rect 4406 54918 4458 54970
rect 4470 54918 4522 54970
rect 34934 54918 34986 54970
rect 34998 54918 35050 54970
rect 35062 54918 35114 54970
rect 35126 54918 35178 54970
rect 35190 54918 35242 54970
rect 45100 54816 45152 54868
rect 41696 54680 41748 54732
rect 42340 54723 42392 54732
rect 42340 54689 42349 54723
rect 42349 54689 42383 54723
rect 42383 54689 42392 54723
rect 42340 54680 42392 54689
rect 43168 54680 43220 54732
rect 1952 54612 2004 54664
rect 43076 54655 43128 54664
rect 43076 54621 43085 54655
rect 43085 54621 43119 54655
rect 43119 54621 43128 54655
rect 43076 54612 43128 54621
rect 42984 54476 43036 54528
rect 43536 54476 43588 54528
rect 19574 54374 19626 54426
rect 19638 54374 19690 54426
rect 19702 54374 19754 54426
rect 19766 54374 19818 54426
rect 19830 54374 19882 54426
rect 50294 54374 50346 54426
rect 50358 54374 50410 54426
rect 50422 54374 50474 54426
rect 50486 54374 50538 54426
rect 50550 54374 50602 54426
rect 1952 54179 2004 54188
rect 1952 54145 1961 54179
rect 1961 54145 1995 54179
rect 1995 54145 2004 54179
rect 1952 54136 2004 54145
rect 46480 54179 46532 54188
rect 2136 54111 2188 54120
rect 2136 54077 2145 54111
rect 2145 54077 2179 54111
rect 2179 54077 2188 54111
rect 2136 54068 2188 54077
rect 2780 54111 2832 54120
rect 2780 54077 2789 54111
rect 2789 54077 2823 54111
rect 2823 54077 2832 54111
rect 2780 54068 2832 54077
rect 46480 54145 46489 54179
rect 46489 54145 46523 54179
rect 46523 54145 46532 54179
rect 46480 54136 46532 54145
rect 47676 54068 47728 54120
rect 46296 53975 46348 53984
rect 46296 53941 46305 53975
rect 46305 53941 46339 53975
rect 46339 53941 46348 53975
rect 46296 53932 46348 53941
rect 4214 53830 4266 53882
rect 4278 53830 4330 53882
rect 4342 53830 4394 53882
rect 4406 53830 4458 53882
rect 4470 53830 4522 53882
rect 34934 53830 34986 53882
rect 34998 53830 35050 53882
rect 35062 53830 35114 53882
rect 35126 53830 35178 53882
rect 35190 53830 35242 53882
rect 2136 53728 2188 53780
rect 46480 53728 46532 53780
rect 49608 53728 49660 53780
rect 45284 53660 45336 53712
rect 2596 53524 2648 53576
rect 42892 53524 42944 53576
rect 45744 53567 45796 53576
rect 45744 53533 45753 53567
rect 45753 53533 45787 53567
rect 45787 53533 45796 53567
rect 45744 53524 45796 53533
rect 45928 53524 45980 53576
rect 47676 53456 47728 53508
rect 45652 53431 45704 53440
rect 45652 53397 45661 53431
rect 45661 53397 45695 53431
rect 45695 53397 45704 53431
rect 45652 53388 45704 53397
rect 19574 53286 19626 53338
rect 19638 53286 19690 53338
rect 19702 53286 19754 53338
rect 19766 53286 19818 53338
rect 19830 53286 19882 53338
rect 50294 53286 50346 53338
rect 50358 53286 50410 53338
rect 50422 53286 50474 53338
rect 50486 53286 50538 53338
rect 50550 53286 50602 53338
rect 44180 53184 44232 53236
rect 46296 53116 46348 53168
rect 49976 53116 50028 53168
rect 42340 53048 42392 53100
rect 42984 53048 43036 53100
rect 48136 53048 48188 53100
rect 48872 53048 48924 53100
rect 42892 53023 42944 53032
rect 42892 52989 42904 53023
rect 42904 52989 42938 53023
rect 42938 52989 42944 53023
rect 42892 52980 42944 52989
rect 43628 52980 43680 53032
rect 46940 52980 46992 53032
rect 47584 52980 47636 53032
rect 47676 52980 47728 53032
rect 47952 52955 48004 52964
rect 47952 52921 47961 52955
rect 47961 52921 47995 52955
rect 47995 52921 48004 52955
rect 47952 52912 48004 52921
rect 49608 52912 49660 52964
rect 45928 52844 45980 52896
rect 47768 52844 47820 52896
rect 49240 52887 49292 52896
rect 49240 52853 49249 52887
rect 49249 52853 49283 52887
rect 49283 52853 49292 52887
rect 50344 53023 50396 53032
rect 50344 52989 50353 53023
rect 50353 52989 50387 53023
rect 50387 52989 50396 53023
rect 50344 52980 50396 52989
rect 49240 52844 49292 52853
rect 50436 52844 50488 52896
rect 51540 52844 51592 52896
rect 4214 52742 4266 52794
rect 4278 52742 4330 52794
rect 4342 52742 4394 52794
rect 4406 52742 4458 52794
rect 4470 52742 4522 52794
rect 34934 52742 34986 52794
rect 34998 52742 35050 52794
rect 35062 52742 35114 52794
rect 35126 52742 35178 52794
rect 35190 52742 35242 52794
rect 42800 52640 42852 52692
rect 43628 52640 43680 52692
rect 42248 52504 42300 52556
rect 46756 52640 46808 52692
rect 46940 52640 46992 52692
rect 48136 52640 48188 52692
rect 48872 52615 48924 52624
rect 48872 52581 48881 52615
rect 48881 52581 48915 52615
rect 48915 52581 48924 52615
rect 48872 52572 48924 52581
rect 50344 52572 50396 52624
rect 42616 52479 42668 52488
rect 42616 52445 42625 52479
rect 42625 52445 42659 52479
rect 42659 52445 42668 52479
rect 42616 52436 42668 52445
rect 45284 52479 45336 52488
rect 45284 52445 45318 52479
rect 45318 52445 45336 52479
rect 45284 52436 45336 52445
rect 46848 52436 46900 52488
rect 47584 52436 47636 52488
rect 47768 52479 47820 52488
rect 47768 52445 47802 52479
rect 47802 52445 47820 52479
rect 47768 52436 47820 52445
rect 49240 52436 49292 52488
rect 49608 52479 49660 52488
rect 49608 52445 49617 52479
rect 49617 52445 49651 52479
rect 49651 52445 49660 52479
rect 49608 52436 49660 52445
rect 49516 52411 49568 52420
rect 49516 52377 49525 52411
rect 49525 52377 49559 52411
rect 49559 52377 49568 52411
rect 50436 52436 50488 52488
rect 49516 52368 49568 52377
rect 49976 52368 50028 52420
rect 42984 52300 43036 52352
rect 43812 52300 43864 52352
rect 50988 52343 51040 52352
rect 50988 52309 50997 52343
rect 50997 52309 51031 52343
rect 51031 52309 51040 52343
rect 50988 52300 51040 52309
rect 19574 52198 19626 52250
rect 19638 52198 19690 52250
rect 19702 52198 19754 52250
rect 19766 52198 19818 52250
rect 19830 52198 19882 52250
rect 50294 52198 50346 52250
rect 50358 52198 50410 52250
rect 50422 52198 50474 52250
rect 50486 52198 50538 52250
rect 50550 52198 50602 52250
rect 42616 52096 42668 52148
rect 43812 52139 43864 52148
rect 43812 52105 43814 52139
rect 43814 52105 43848 52139
rect 43848 52105 43864 52139
rect 43812 52096 43864 52105
rect 45652 52096 45704 52148
rect 45744 52096 45796 52148
rect 46020 52096 46072 52148
rect 47952 52139 48004 52148
rect 47952 52105 47961 52139
rect 47961 52105 47995 52139
rect 47995 52105 48004 52139
rect 47952 52096 48004 52105
rect 49516 52139 49568 52148
rect 49516 52105 49525 52139
rect 49525 52105 49559 52139
rect 49559 52105 49568 52139
rect 49516 52096 49568 52105
rect 48320 52028 48372 52080
rect 48872 52028 48924 52080
rect 49240 52028 49292 52080
rect 42800 51960 42852 52012
rect 43536 51935 43588 51944
rect 43536 51901 43545 51935
rect 43545 51901 43579 51935
rect 43579 51901 43588 51935
rect 43536 51892 43588 51901
rect 45928 51960 45980 52012
rect 46664 51960 46716 52012
rect 46940 52003 46992 52012
rect 46940 51969 46949 52003
rect 46949 51969 46983 52003
rect 46983 51969 46992 52003
rect 46940 51960 46992 51969
rect 49608 51960 49660 52012
rect 51540 52003 51592 52012
rect 51540 51969 51549 52003
rect 51549 51969 51583 52003
rect 51583 51969 51592 52003
rect 51540 51960 51592 51969
rect 42340 51756 42392 51808
rect 46112 51892 46164 51944
rect 49976 51867 50028 51876
rect 49976 51833 49985 51867
rect 49985 51833 50019 51867
rect 50019 51833 50028 51867
rect 49976 51824 50028 51833
rect 46664 51799 46716 51808
rect 46664 51765 46673 51799
rect 46673 51765 46707 51799
rect 46707 51765 46716 51799
rect 46664 51756 46716 51765
rect 46848 51756 46900 51808
rect 49424 51756 49476 51808
rect 50620 51756 50672 51808
rect 52920 51756 52972 51808
rect 4214 51654 4266 51706
rect 4278 51654 4330 51706
rect 4342 51654 4394 51706
rect 4406 51654 4458 51706
rect 4470 51654 4522 51706
rect 34934 51654 34986 51706
rect 34998 51654 35050 51706
rect 35062 51654 35114 51706
rect 35126 51654 35178 51706
rect 35190 51654 35242 51706
rect 46112 51552 46164 51604
rect 44732 51348 44784 51400
rect 45836 51416 45888 51468
rect 45652 51348 45704 51400
rect 45928 51348 45980 51400
rect 46848 51348 46900 51400
rect 48596 51348 48648 51400
rect 50988 51348 51040 51400
rect 48320 51280 48372 51332
rect 45468 51212 45520 51264
rect 50804 51255 50856 51264
rect 50804 51221 50813 51255
rect 50813 51221 50847 51255
rect 50847 51221 50856 51255
rect 50804 51212 50856 51221
rect 19574 51110 19626 51162
rect 19638 51110 19690 51162
rect 19702 51110 19754 51162
rect 19766 51110 19818 51162
rect 19830 51110 19882 51162
rect 50294 51110 50346 51162
rect 50358 51110 50410 51162
rect 50422 51110 50474 51162
rect 50486 51110 50538 51162
rect 50550 51110 50602 51162
rect 49976 51008 50028 51060
rect 44732 50915 44784 50924
rect 44732 50881 44741 50915
rect 44741 50881 44775 50915
rect 44775 50881 44784 50915
rect 44732 50872 44784 50881
rect 46112 50940 46164 50992
rect 45836 50915 45888 50924
rect 45836 50881 45845 50915
rect 45845 50881 45879 50915
rect 45879 50881 45888 50915
rect 45836 50872 45888 50881
rect 46020 50915 46072 50924
rect 46020 50881 46029 50915
rect 46029 50881 46063 50915
rect 46063 50881 46072 50915
rect 46020 50872 46072 50881
rect 48596 50872 48648 50924
rect 49424 50915 49476 50924
rect 49424 50881 49433 50915
rect 49433 50881 49467 50915
rect 49467 50881 49476 50915
rect 49424 50872 49476 50881
rect 50620 50872 50672 50924
rect 43812 50668 43864 50720
rect 46020 50711 46072 50720
rect 46020 50677 46029 50711
rect 46029 50677 46063 50711
rect 46063 50677 46072 50711
rect 46020 50668 46072 50677
rect 49240 50711 49292 50720
rect 49240 50677 49249 50711
rect 49249 50677 49283 50711
rect 49283 50677 49292 50711
rect 49240 50668 49292 50677
rect 50620 50668 50672 50720
rect 4214 50566 4266 50618
rect 4278 50566 4330 50618
rect 4342 50566 4394 50618
rect 4406 50566 4458 50618
rect 4470 50566 4522 50618
rect 34934 50566 34986 50618
rect 34998 50566 35050 50618
rect 35062 50566 35114 50618
rect 35126 50566 35178 50618
rect 35190 50566 35242 50618
rect 49976 50396 50028 50448
rect 36268 50260 36320 50312
rect 40500 50260 40552 50312
rect 47676 50303 47728 50312
rect 47676 50269 47685 50303
rect 47685 50269 47719 50303
rect 47719 50269 47728 50303
rect 47676 50260 47728 50269
rect 48136 50303 48188 50312
rect 48136 50269 48145 50303
rect 48145 50269 48179 50303
rect 48179 50269 48188 50303
rect 48136 50260 48188 50269
rect 37924 50192 37976 50244
rect 48044 50192 48096 50244
rect 39488 50124 39540 50176
rect 47492 50167 47544 50176
rect 47492 50133 47501 50167
rect 47501 50133 47535 50167
rect 47535 50133 47544 50167
rect 47492 50124 47544 50133
rect 19574 50022 19626 50074
rect 19638 50022 19690 50074
rect 19702 50022 19754 50074
rect 19766 50022 19818 50074
rect 19830 50022 19882 50074
rect 50294 50022 50346 50074
rect 50358 50022 50410 50074
rect 50422 50022 50474 50074
rect 50486 50022 50538 50074
rect 50550 50022 50602 50074
rect 37924 49963 37976 49972
rect 37924 49929 37933 49963
rect 37933 49929 37967 49963
rect 37967 49929 37976 49963
rect 37924 49920 37976 49929
rect 43720 49963 43772 49972
rect 43720 49929 43735 49963
rect 43735 49929 43769 49963
rect 43769 49929 43772 49963
rect 43720 49920 43772 49929
rect 50712 49920 50764 49972
rect 53196 49920 53248 49972
rect 47492 49852 47544 49904
rect 38108 49827 38160 49836
rect 38108 49793 38117 49827
rect 38117 49793 38151 49827
rect 38151 49793 38160 49827
rect 38108 49784 38160 49793
rect 39488 49827 39540 49836
rect 1952 49759 2004 49768
rect 1952 49725 1961 49759
rect 1961 49725 1995 49759
rect 1995 49725 2004 49759
rect 1952 49716 2004 49725
rect 2136 49759 2188 49768
rect 2136 49725 2145 49759
rect 2145 49725 2179 49759
rect 2179 49725 2188 49759
rect 2136 49716 2188 49725
rect 2780 49759 2832 49768
rect 2780 49725 2789 49759
rect 2789 49725 2823 49759
rect 2823 49725 2832 49759
rect 2780 49716 2832 49725
rect 37556 49716 37608 49768
rect 39488 49793 39497 49827
rect 39497 49793 39531 49827
rect 39531 49793 39540 49827
rect 39488 49784 39540 49793
rect 40500 49827 40552 49836
rect 40500 49793 40509 49827
rect 40509 49793 40543 49827
rect 40543 49793 40552 49827
rect 40500 49784 40552 49793
rect 40776 49827 40828 49836
rect 40776 49793 40810 49827
rect 40810 49793 40828 49827
rect 40776 49784 40828 49793
rect 42340 49784 42392 49836
rect 43812 49716 43864 49768
rect 44180 49716 44232 49768
rect 47584 49759 47636 49768
rect 47584 49725 47593 49759
rect 47593 49725 47627 49759
rect 47627 49725 47636 49759
rect 47584 49716 47636 49725
rect 50160 49716 50212 49768
rect 50804 49759 50856 49768
rect 50804 49725 50816 49759
rect 50816 49725 50850 49759
rect 50850 49725 50856 49759
rect 51080 49759 51132 49768
rect 50804 49716 50856 49725
rect 51080 49725 51089 49759
rect 51089 49725 51123 49759
rect 51123 49725 51132 49759
rect 51080 49716 51132 49725
rect 38568 49648 38620 49700
rect 39856 49580 39908 49632
rect 41420 49580 41472 49632
rect 42708 49580 42760 49632
rect 45100 49623 45152 49632
rect 45100 49589 45109 49623
rect 45109 49589 45143 49623
rect 45143 49589 45152 49623
rect 45100 49580 45152 49589
rect 48596 49580 48648 49632
rect 4214 49478 4266 49530
rect 4278 49478 4330 49530
rect 4342 49478 4394 49530
rect 4406 49478 4458 49530
rect 4470 49478 4522 49530
rect 34934 49478 34986 49530
rect 34998 49478 35050 49530
rect 35062 49478 35114 49530
rect 35126 49478 35178 49530
rect 35190 49478 35242 49530
rect 1952 49376 2004 49428
rect 39488 49376 39540 49428
rect 36268 49283 36320 49292
rect 36268 49249 36277 49283
rect 36277 49249 36311 49283
rect 36311 49249 36320 49283
rect 36268 49240 36320 49249
rect 40224 49308 40276 49360
rect 50160 49376 50212 49428
rect 50804 49376 50856 49428
rect 51080 49376 51132 49428
rect 45468 49283 45520 49292
rect 45468 49249 45480 49283
rect 45480 49249 45514 49283
rect 45514 49249 45520 49283
rect 45468 49240 45520 49249
rect 48136 49240 48188 49292
rect 39856 49172 39908 49224
rect 40316 49215 40368 49224
rect 40316 49181 40325 49215
rect 40325 49181 40359 49215
rect 40359 49181 40368 49215
rect 40868 49215 40920 49224
rect 40316 49172 40368 49181
rect 36728 49104 36780 49156
rect 39396 49104 39448 49156
rect 39488 49104 39540 49156
rect 40132 49104 40184 49156
rect 40868 49181 40877 49215
rect 40877 49181 40911 49215
rect 40911 49181 40920 49215
rect 40868 49172 40920 49181
rect 41420 49172 41472 49224
rect 41604 49215 41656 49224
rect 41604 49181 41613 49215
rect 41613 49181 41647 49215
rect 41647 49181 41656 49215
rect 41604 49172 41656 49181
rect 42340 49172 42392 49224
rect 45008 49215 45060 49224
rect 45008 49181 45017 49215
rect 45017 49181 45051 49215
rect 45051 49181 45060 49215
rect 45008 49172 45060 49181
rect 45100 49172 45152 49224
rect 47768 49215 47820 49224
rect 47768 49181 47777 49215
rect 47777 49181 47811 49215
rect 47811 49181 47820 49215
rect 50160 49215 50212 49224
rect 47768 49172 47820 49181
rect 50160 49181 50169 49215
rect 50169 49181 50203 49215
rect 50203 49181 50212 49215
rect 50160 49172 50212 49181
rect 50620 49283 50672 49292
rect 50620 49249 50632 49283
rect 50632 49249 50666 49283
rect 50666 49249 50672 49283
rect 50620 49240 50672 49249
rect 52644 49240 52696 49292
rect 52920 49283 52972 49292
rect 52920 49249 52932 49283
rect 52932 49249 52966 49283
rect 52966 49249 52972 49283
rect 53196 49283 53248 49292
rect 52920 49240 52972 49249
rect 53196 49249 53205 49283
rect 53205 49249 53239 49283
rect 53239 49249 53248 49283
rect 53196 49240 53248 49249
rect 51172 49172 51224 49224
rect 37924 49036 37976 49088
rect 40500 49036 40552 49088
rect 41328 49079 41380 49088
rect 41328 49045 41343 49079
rect 41343 49045 41377 49079
rect 41377 49045 41380 49079
rect 41328 49036 41380 49045
rect 43168 49036 43220 49088
rect 46204 49036 46256 49088
rect 46848 49079 46900 49088
rect 46848 49045 46857 49079
rect 46857 49045 46891 49079
rect 46891 49045 46900 49079
rect 46848 49036 46900 49045
rect 48964 49036 49016 49088
rect 49608 49079 49660 49088
rect 49608 49045 49617 49079
rect 49617 49045 49651 49079
rect 49651 49045 49660 49079
rect 49608 49036 49660 49045
rect 50620 49079 50672 49088
rect 50620 49045 50635 49079
rect 50635 49045 50669 49079
rect 50669 49045 50672 49079
rect 50620 49036 50672 49045
rect 50804 49036 50856 49088
rect 52276 49036 52328 49088
rect 19574 48934 19626 48986
rect 19638 48934 19690 48986
rect 19702 48934 19754 48986
rect 19766 48934 19818 48986
rect 19830 48934 19882 48986
rect 50294 48934 50346 48986
rect 50358 48934 50410 48986
rect 50422 48934 50474 48986
rect 50486 48934 50538 48986
rect 50550 48934 50602 48986
rect 2136 48832 2188 48884
rect 36728 48875 36780 48884
rect 36728 48841 36737 48875
rect 36737 48841 36771 48875
rect 36771 48841 36780 48875
rect 36728 48832 36780 48841
rect 37556 48875 37608 48884
rect 37556 48841 37565 48875
rect 37565 48841 37599 48875
rect 37599 48841 37608 48875
rect 37556 48832 37608 48841
rect 38108 48832 38160 48884
rect 39396 48875 39448 48884
rect 39396 48841 39405 48875
rect 39405 48841 39439 48875
rect 39439 48841 39448 48875
rect 39396 48832 39448 48841
rect 39672 48832 39724 48884
rect 40776 48832 40828 48884
rect 41052 48832 41104 48884
rect 41328 48832 41380 48884
rect 43628 48832 43680 48884
rect 44180 48832 44232 48884
rect 47584 48832 47636 48884
rect 48964 48832 49016 48884
rect 2504 48739 2556 48748
rect 2504 48705 2513 48739
rect 2513 48705 2547 48739
rect 2547 48705 2556 48739
rect 2504 48696 2556 48705
rect 37924 48807 37976 48816
rect 37924 48773 37933 48807
rect 37933 48773 37967 48807
rect 37967 48773 37976 48807
rect 37924 48764 37976 48773
rect 38568 48764 38620 48816
rect 37832 48696 37884 48748
rect 40224 48764 40276 48816
rect 48596 48764 48648 48816
rect 51172 48832 51224 48884
rect 50620 48764 50672 48816
rect 52644 48764 52696 48816
rect 39488 48696 39540 48748
rect 40316 48696 40368 48748
rect 40500 48739 40552 48748
rect 40500 48705 40509 48739
rect 40509 48705 40543 48739
rect 40543 48705 40552 48739
rect 40500 48696 40552 48705
rect 40868 48696 40920 48748
rect 42340 48696 42392 48748
rect 43168 48739 43220 48748
rect 43168 48705 43177 48739
rect 43177 48705 43211 48739
rect 43211 48705 43220 48739
rect 43168 48696 43220 48705
rect 45100 48696 45152 48748
rect 36452 48671 36504 48680
rect 36452 48637 36461 48671
rect 36461 48637 36495 48671
rect 36495 48637 36504 48671
rect 36452 48628 36504 48637
rect 37464 48560 37516 48612
rect 38844 48671 38896 48680
rect 38844 48637 38853 48671
rect 38853 48637 38887 48671
rect 38887 48637 38896 48671
rect 38844 48628 38896 48637
rect 39948 48671 40000 48680
rect 39948 48637 39957 48671
rect 39957 48637 39991 48671
rect 39991 48637 40000 48671
rect 39948 48628 40000 48637
rect 39856 48560 39908 48612
rect 42892 48671 42944 48680
rect 42892 48637 42904 48671
rect 42904 48637 42938 48671
rect 42938 48637 42944 48671
rect 44732 48671 44784 48680
rect 42892 48628 42944 48637
rect 44732 48637 44741 48671
rect 44741 48637 44775 48671
rect 44775 48637 44784 48671
rect 44732 48628 44784 48637
rect 47768 48628 47820 48680
rect 49240 48628 49292 48680
rect 49332 48671 49384 48680
rect 49332 48637 49341 48671
rect 49341 48637 49375 48671
rect 49375 48637 49384 48671
rect 49332 48628 49384 48637
rect 48044 48603 48096 48612
rect 48044 48569 48053 48603
rect 48053 48569 48087 48603
rect 48087 48569 48096 48603
rect 48044 48560 48096 48569
rect 37556 48492 37608 48544
rect 39488 48492 39540 48544
rect 48412 48492 48464 48544
rect 4214 48390 4266 48442
rect 4278 48390 4330 48442
rect 4342 48390 4394 48442
rect 4406 48390 4458 48442
rect 4470 48390 4522 48442
rect 34934 48390 34986 48442
rect 34998 48390 35050 48442
rect 35062 48390 35114 48442
rect 35126 48390 35178 48442
rect 35190 48390 35242 48442
rect 37464 48331 37516 48340
rect 37464 48297 37473 48331
rect 37473 48297 37507 48331
rect 37507 48297 37516 48331
rect 37464 48288 37516 48297
rect 45008 48288 45060 48340
rect 40224 48152 40276 48204
rect 47768 48288 47820 48340
rect 48136 48288 48188 48340
rect 49332 48220 49384 48272
rect 46020 48152 46072 48204
rect 46388 48152 46440 48204
rect 46848 48152 46900 48204
rect 1952 48084 2004 48136
rect 36728 48084 36780 48136
rect 37832 48084 37884 48136
rect 39304 48084 39356 48136
rect 39948 48084 40000 48136
rect 48412 48127 48464 48136
rect 48412 48093 48421 48127
rect 48421 48093 48455 48127
rect 48455 48093 48464 48127
rect 48412 48084 48464 48093
rect 38568 48016 38620 48068
rect 37372 47948 37424 48000
rect 46204 47991 46256 48000
rect 46204 47957 46219 47991
rect 46219 47957 46253 47991
rect 46253 47957 46256 47991
rect 46204 47948 46256 47957
rect 19574 47846 19626 47898
rect 19638 47846 19690 47898
rect 19702 47846 19754 47898
rect 19766 47846 19818 47898
rect 19830 47846 19882 47898
rect 50294 47846 50346 47898
rect 50358 47846 50410 47898
rect 50422 47846 50474 47898
rect 50486 47846 50538 47898
rect 50550 47846 50602 47898
rect 40316 47744 40368 47796
rect 41052 47744 41104 47796
rect 41604 47744 41656 47796
rect 47676 47744 47728 47796
rect 44732 47676 44784 47728
rect 1952 47651 2004 47660
rect 1952 47617 1961 47651
rect 1961 47617 1995 47651
rect 1995 47617 2004 47651
rect 1952 47608 2004 47617
rect 36452 47608 36504 47660
rect 36728 47651 36780 47660
rect 36728 47617 36737 47651
rect 36737 47617 36771 47651
rect 36771 47617 36780 47651
rect 36728 47608 36780 47617
rect 37372 47608 37424 47660
rect 38568 47608 38620 47660
rect 46388 47651 46440 47660
rect 2412 47540 2464 47592
rect 2780 47583 2832 47592
rect 2780 47549 2789 47583
rect 2789 47549 2823 47583
rect 2823 47549 2832 47583
rect 2780 47540 2832 47549
rect 37556 47540 37608 47592
rect 38476 47540 38528 47592
rect 40224 47540 40276 47592
rect 46388 47617 46397 47651
rect 46397 47617 46431 47651
rect 46431 47617 46440 47651
rect 46388 47608 46440 47617
rect 50804 47608 50856 47660
rect 41880 47540 41932 47592
rect 36360 47447 36412 47456
rect 36360 47413 36369 47447
rect 36369 47413 36403 47447
rect 36403 47413 36412 47447
rect 36360 47404 36412 47413
rect 38200 47404 38252 47456
rect 4214 47302 4266 47354
rect 4278 47302 4330 47354
rect 4342 47302 4394 47354
rect 4406 47302 4458 47354
rect 4470 47302 4522 47354
rect 34934 47302 34986 47354
rect 34998 47302 35050 47354
rect 35062 47302 35114 47354
rect 35126 47302 35178 47354
rect 35190 47302 35242 47354
rect 2412 47243 2464 47252
rect 2412 47209 2421 47243
rect 2421 47209 2455 47243
rect 2455 47209 2464 47243
rect 2412 47200 2464 47209
rect 38200 47243 38252 47252
rect 38200 47209 38209 47243
rect 38209 47209 38243 47243
rect 38243 47209 38252 47243
rect 38200 47200 38252 47209
rect 39304 47243 39356 47252
rect 39304 47209 39313 47243
rect 39313 47209 39347 47243
rect 39347 47209 39356 47243
rect 39304 47200 39356 47209
rect 36360 47132 36412 47184
rect 2596 46996 2648 47048
rect 8852 46996 8904 47048
rect 36268 46996 36320 47048
rect 37648 46996 37700 47048
rect 40132 47107 40184 47116
rect 40132 47073 40141 47107
rect 40141 47073 40175 47107
rect 40175 47073 40184 47107
rect 40132 47064 40184 47073
rect 42800 47064 42852 47116
rect 44732 47200 44784 47252
rect 52736 47200 52788 47252
rect 50804 47107 50856 47116
rect 50804 47073 50813 47107
rect 50813 47073 50847 47107
rect 50847 47073 50856 47107
rect 50804 47064 50856 47073
rect 52276 47107 52328 47116
rect 52276 47073 52285 47107
rect 52285 47073 52319 47107
rect 52319 47073 52328 47107
rect 52276 47064 52328 47073
rect 52644 47064 52696 47116
rect 52920 47064 52972 47116
rect 38476 47039 38528 47048
rect 38476 47005 38485 47039
rect 38485 47005 38519 47039
rect 38519 47005 38528 47039
rect 39120 47039 39172 47048
rect 38476 46996 38528 47005
rect 39120 47005 39129 47039
rect 39129 47005 39163 47039
rect 39163 47005 39172 47039
rect 39120 46996 39172 47005
rect 39672 46996 39724 47048
rect 43076 46996 43128 47048
rect 43628 46996 43680 47048
rect 44364 46996 44416 47048
rect 51080 47039 51132 47048
rect 51080 47005 51089 47039
rect 51089 47005 51123 47039
rect 51123 47005 51132 47039
rect 58164 47039 58216 47048
rect 51080 46996 51132 47005
rect 44456 46903 44508 46912
rect 44456 46869 44465 46903
rect 44465 46869 44499 46903
rect 44499 46869 44508 46903
rect 44456 46860 44508 46869
rect 58164 47005 58173 47039
rect 58173 47005 58207 47039
rect 58207 47005 58216 47039
rect 58164 46996 58216 47005
rect 19574 46758 19626 46810
rect 19638 46758 19690 46810
rect 19702 46758 19754 46810
rect 19766 46758 19818 46810
rect 19830 46758 19882 46810
rect 50294 46758 50346 46810
rect 50358 46758 50410 46810
rect 50422 46758 50474 46810
rect 50486 46758 50538 46810
rect 50550 46758 50602 46810
rect 40316 46656 40368 46708
rect 41880 46699 41932 46708
rect 37648 46588 37700 46640
rect 38660 46520 38712 46572
rect 39120 46520 39172 46572
rect 41880 46665 41889 46699
rect 41889 46665 41923 46699
rect 41923 46665 41932 46699
rect 41880 46656 41932 46665
rect 44364 46656 44416 46708
rect 46204 46656 46256 46708
rect 48044 46656 48096 46708
rect 49424 46656 49476 46708
rect 46204 46520 46256 46572
rect 49608 46520 49660 46572
rect 53012 46588 53064 46640
rect 37372 46384 37424 46436
rect 37464 46316 37516 46368
rect 39856 46316 39908 46368
rect 41788 46452 41840 46504
rect 42340 46452 42392 46504
rect 43076 46495 43128 46504
rect 43076 46461 43088 46495
rect 43088 46461 43122 46495
rect 43122 46461 43128 46495
rect 43076 46452 43128 46461
rect 40224 46316 40276 46368
rect 47032 46452 47084 46504
rect 44180 46384 44232 46436
rect 47768 46316 47820 46368
rect 50804 46384 50856 46436
rect 53288 46427 53340 46436
rect 53288 46393 53297 46427
rect 53297 46393 53331 46427
rect 53331 46393 53340 46427
rect 53288 46384 53340 46393
rect 50620 46316 50672 46368
rect 52736 46316 52788 46368
rect 4214 46214 4266 46266
rect 4278 46214 4330 46266
rect 4342 46214 4394 46266
rect 4406 46214 4458 46266
rect 4470 46214 4522 46266
rect 34934 46214 34986 46266
rect 34998 46214 35050 46266
rect 35062 46214 35114 46266
rect 35126 46214 35178 46266
rect 35190 46214 35242 46266
rect 53288 46044 53340 46096
rect 36268 46019 36320 46028
rect 36268 45985 36277 46019
rect 36277 45985 36311 46019
rect 36311 45985 36320 46019
rect 36268 45976 36320 45985
rect 38660 45976 38712 46028
rect 40132 45976 40184 46028
rect 44732 45976 44784 46028
rect 47768 46019 47820 46028
rect 47768 45985 47777 46019
rect 47777 45985 47811 46019
rect 47811 45985 47820 46019
rect 47768 45976 47820 45985
rect 48044 45976 48096 46028
rect 48228 46019 48280 46028
rect 48228 45985 48240 46019
rect 48240 45985 48274 46019
rect 48274 45985 48280 46019
rect 48228 45976 48280 45985
rect 50988 45976 51040 46028
rect 52920 45976 52972 46028
rect 53196 45976 53248 46028
rect 36360 45908 36412 45960
rect 44180 45951 44232 45960
rect 44180 45917 44189 45951
rect 44189 45917 44223 45951
rect 44223 45917 44232 45951
rect 44180 45908 44232 45917
rect 37280 45840 37332 45892
rect 50896 45908 50948 45960
rect 52736 45951 52788 45960
rect 37648 45815 37700 45824
rect 37648 45781 37657 45815
rect 37657 45781 37691 45815
rect 37691 45781 37700 45815
rect 37648 45772 37700 45781
rect 43076 45772 43128 45824
rect 45928 45883 45980 45892
rect 45928 45849 45962 45883
rect 45962 45849 45980 45883
rect 45928 45840 45980 45849
rect 49240 45840 49292 45892
rect 52736 45917 52745 45951
rect 52745 45917 52779 45951
rect 52779 45917 52788 45951
rect 52736 45908 52788 45917
rect 47124 45772 47176 45824
rect 48044 45772 48096 45824
rect 49884 45772 49936 45824
rect 19574 45670 19626 45722
rect 19638 45670 19690 45722
rect 19702 45670 19754 45722
rect 19766 45670 19818 45722
rect 19830 45670 19882 45722
rect 50294 45670 50346 45722
rect 50358 45670 50410 45722
rect 50422 45670 50474 45722
rect 50486 45670 50538 45722
rect 50550 45670 50602 45722
rect 40316 45568 40368 45620
rect 41788 45611 41840 45620
rect 41788 45577 41797 45611
rect 41797 45577 41831 45611
rect 41831 45577 41840 45611
rect 41788 45568 41840 45577
rect 49240 45568 49292 45620
rect 49424 45568 49476 45620
rect 52736 45611 52788 45620
rect 52736 45577 52745 45611
rect 52745 45577 52779 45611
rect 52779 45577 52788 45611
rect 52736 45568 52788 45577
rect 53288 45568 53340 45620
rect 37280 45543 37332 45552
rect 37280 45509 37289 45543
rect 37289 45509 37323 45543
rect 37323 45509 37332 45543
rect 37280 45500 37332 45509
rect 47032 45500 47084 45552
rect 37464 45475 37516 45484
rect 37464 45441 37473 45475
rect 37473 45441 37507 45475
rect 37507 45441 37516 45475
rect 37464 45432 37516 45441
rect 37648 45432 37700 45484
rect 44180 45432 44232 45484
rect 44456 45432 44508 45484
rect 45560 45475 45612 45484
rect 45560 45441 45569 45475
rect 45569 45441 45603 45475
rect 45603 45441 45612 45475
rect 45560 45432 45612 45441
rect 39856 45364 39908 45416
rect 41696 45364 41748 45416
rect 45468 45407 45520 45416
rect 45468 45373 45477 45407
rect 45477 45373 45511 45407
rect 45511 45373 45520 45407
rect 45468 45364 45520 45373
rect 47400 45432 47452 45484
rect 52828 45432 52880 45484
rect 47124 45364 47176 45416
rect 50620 45364 50672 45416
rect 50804 45407 50856 45416
rect 50804 45373 50813 45407
rect 50813 45373 50847 45407
rect 50847 45373 50856 45407
rect 50804 45364 50856 45373
rect 51080 45364 51132 45416
rect 1952 45228 2004 45280
rect 37372 45228 37424 45280
rect 43904 45271 43956 45280
rect 43904 45237 43913 45271
rect 43913 45237 43947 45271
rect 43947 45237 43956 45271
rect 43904 45228 43956 45237
rect 44456 45228 44508 45280
rect 46664 45228 46716 45280
rect 46756 45271 46808 45280
rect 46756 45237 46765 45271
rect 46765 45237 46799 45271
rect 46799 45237 46808 45271
rect 46756 45228 46808 45237
rect 53012 45228 53064 45280
rect 4214 45126 4266 45178
rect 4278 45126 4330 45178
rect 4342 45126 4394 45178
rect 4406 45126 4458 45178
rect 4470 45126 4522 45178
rect 34934 45126 34986 45178
rect 34998 45126 35050 45178
rect 35062 45126 35114 45178
rect 35126 45126 35178 45178
rect 35190 45126 35242 45178
rect 41696 45067 41748 45076
rect 41696 45033 41705 45067
rect 41705 45033 41739 45067
rect 41739 45033 41748 45067
rect 41696 45024 41748 45033
rect 45928 45024 45980 45076
rect 46664 45024 46716 45076
rect 47400 45067 47452 45076
rect 47400 45033 47409 45067
rect 47409 45033 47443 45067
rect 47443 45033 47452 45067
rect 47400 45024 47452 45033
rect 36452 44888 36504 44940
rect 39488 44888 39540 44940
rect 45468 44888 45520 44940
rect 2504 44863 2556 44872
rect 2504 44829 2513 44863
rect 2513 44829 2547 44863
rect 2547 44829 2556 44863
rect 2504 44820 2556 44829
rect 37372 44820 37424 44872
rect 37464 44863 37516 44872
rect 37464 44829 37473 44863
rect 37473 44829 37507 44863
rect 37507 44829 37516 44863
rect 37464 44820 37516 44829
rect 39856 44863 39908 44872
rect 39856 44829 39865 44863
rect 39865 44829 39899 44863
rect 39899 44829 39908 44863
rect 39856 44820 39908 44829
rect 41696 44820 41748 44872
rect 43076 44863 43128 44872
rect 43076 44829 43085 44863
rect 43085 44829 43119 44863
rect 43119 44829 43128 44863
rect 43076 44820 43128 44829
rect 45560 44820 45612 44872
rect 46296 44863 46348 44872
rect 46296 44829 46305 44863
rect 46305 44829 46339 44863
rect 46339 44829 46348 44863
rect 46296 44820 46348 44829
rect 46940 44888 46992 44940
rect 50160 44888 50212 44940
rect 50896 45024 50948 45076
rect 46572 44863 46624 44872
rect 46572 44829 46581 44863
rect 46581 44829 46615 44863
rect 46615 44829 46624 44863
rect 46572 44820 46624 44829
rect 46848 44820 46900 44872
rect 47676 44863 47728 44872
rect 47676 44829 47685 44863
rect 47685 44829 47719 44863
rect 47719 44829 47728 44863
rect 48044 44863 48096 44872
rect 47676 44820 47728 44829
rect 48044 44829 48053 44863
rect 48053 44829 48087 44863
rect 48087 44829 48096 44863
rect 48044 44820 48096 44829
rect 49884 44820 49936 44872
rect 43720 44752 43772 44804
rect 47124 44752 47176 44804
rect 52368 44752 52420 44804
rect 2136 44684 2188 44736
rect 37004 44727 37056 44736
rect 37004 44693 37013 44727
rect 37013 44693 37047 44727
rect 37047 44693 37056 44727
rect 37004 44684 37056 44693
rect 38660 44684 38712 44736
rect 40316 44727 40368 44736
rect 40316 44693 40331 44727
rect 40331 44693 40365 44727
rect 40365 44693 40368 44727
rect 44456 44727 44508 44736
rect 40316 44684 40368 44693
rect 44456 44693 44465 44727
rect 44465 44693 44499 44727
rect 44499 44693 44508 44727
rect 44456 44684 44508 44693
rect 51448 44727 51500 44736
rect 51448 44693 51457 44727
rect 51457 44693 51491 44727
rect 51491 44693 51500 44727
rect 51448 44684 51500 44693
rect 52736 44684 52788 44736
rect 19574 44582 19626 44634
rect 19638 44582 19690 44634
rect 19702 44582 19754 44634
rect 19766 44582 19818 44634
rect 19830 44582 19882 44634
rect 50294 44582 50346 44634
rect 50358 44582 50410 44634
rect 50422 44582 50474 44634
rect 50486 44582 50538 44634
rect 50550 44582 50602 44634
rect 39488 44523 39540 44532
rect 39488 44489 39513 44523
rect 39513 44489 39540 44523
rect 39672 44523 39724 44532
rect 39488 44480 39540 44489
rect 39672 44489 39681 44523
rect 39681 44489 39715 44523
rect 39715 44489 39724 44523
rect 39672 44480 39724 44489
rect 40132 44523 40184 44532
rect 40132 44489 40141 44523
rect 40141 44489 40175 44523
rect 40175 44489 40184 44523
rect 40132 44480 40184 44489
rect 43720 44523 43772 44532
rect 43720 44489 43729 44523
rect 43729 44489 43763 44523
rect 43763 44489 43772 44523
rect 43720 44480 43772 44489
rect 49424 44480 49476 44532
rect 53012 44523 53064 44532
rect 53012 44489 53021 44523
rect 53021 44489 53055 44523
rect 53055 44489 53064 44523
rect 53012 44480 53064 44489
rect 2136 44455 2188 44464
rect 2136 44421 2145 44455
rect 2145 44421 2179 44455
rect 2179 44421 2188 44455
rect 2136 44412 2188 44421
rect 37004 44412 37056 44464
rect 1952 44387 2004 44396
rect 1952 44353 1961 44387
rect 1961 44353 1995 44387
rect 1995 44353 2004 44387
rect 1952 44344 2004 44353
rect 36268 44344 36320 44396
rect 37280 44387 37332 44396
rect 37280 44353 37289 44387
rect 37289 44353 37323 44387
rect 37323 44353 37332 44387
rect 37280 44344 37332 44353
rect 38660 44344 38712 44396
rect 41696 44344 41748 44396
rect 43904 44387 43956 44396
rect 43904 44353 43913 44387
rect 43913 44353 43947 44387
rect 43947 44353 43956 44387
rect 43904 44344 43956 44353
rect 44456 44344 44508 44396
rect 45376 44344 45428 44396
rect 46940 44412 46992 44464
rect 52736 44455 52788 44464
rect 52736 44421 52745 44455
rect 52745 44421 52779 44455
rect 52779 44421 52788 44455
rect 52736 44412 52788 44421
rect 46296 44387 46348 44396
rect 46296 44353 46305 44387
rect 46305 44353 46339 44387
rect 46339 44353 46348 44387
rect 46296 44344 46348 44353
rect 2780 44319 2832 44328
rect 2780 44285 2789 44319
rect 2789 44285 2823 44319
rect 2823 44285 2832 44319
rect 2780 44276 2832 44285
rect 41512 44276 41564 44328
rect 42708 44276 42760 44328
rect 44180 44276 44232 44328
rect 46848 44344 46900 44396
rect 49884 44387 49936 44396
rect 49884 44353 49893 44387
rect 49893 44353 49927 44387
rect 49927 44353 49936 44387
rect 49884 44344 49936 44353
rect 53012 44387 53064 44396
rect 53012 44353 53021 44387
rect 53021 44353 53055 44387
rect 53055 44353 53064 44387
rect 53012 44344 53064 44353
rect 45284 44208 45336 44260
rect 46756 44208 46808 44260
rect 39488 44183 39540 44192
rect 39488 44149 39497 44183
rect 39497 44149 39531 44183
rect 39531 44149 39540 44183
rect 39488 44140 39540 44149
rect 49700 44276 49752 44328
rect 50620 44276 50672 44328
rect 51448 44276 51500 44328
rect 50068 44140 50120 44192
rect 50804 44140 50856 44192
rect 52368 44140 52420 44192
rect 4214 44038 4266 44090
rect 4278 44038 4330 44090
rect 4342 44038 4394 44090
rect 4406 44038 4458 44090
rect 4470 44038 4522 44090
rect 34934 44038 34986 44090
rect 34998 44038 35050 44090
rect 35062 44038 35114 44090
rect 35126 44038 35178 44090
rect 35190 44038 35242 44090
rect 37280 43936 37332 43988
rect 46572 43936 46624 43988
rect 36452 43868 36504 43920
rect 37924 43868 37976 43920
rect 41512 43843 41564 43852
rect 41512 43809 41521 43843
rect 41521 43809 41555 43843
rect 41555 43809 41564 43843
rect 41512 43800 41564 43809
rect 37464 43775 37516 43784
rect 37464 43741 37473 43775
rect 37473 43741 37507 43775
rect 37507 43741 37516 43775
rect 37464 43732 37516 43741
rect 36912 43596 36964 43648
rect 37648 43732 37700 43784
rect 38292 43775 38344 43784
rect 38292 43741 38301 43775
rect 38301 43741 38335 43775
rect 38335 43741 38344 43775
rect 38292 43732 38344 43741
rect 39488 43732 39540 43784
rect 40500 43732 40552 43784
rect 44180 43732 44232 43784
rect 45284 43732 45336 43784
rect 47032 43732 47084 43784
rect 47676 43732 47728 43784
rect 37924 43664 37976 43716
rect 38660 43596 38712 43648
rect 44272 43639 44324 43648
rect 44272 43605 44281 43639
rect 44281 43605 44315 43639
rect 44315 43605 44324 43639
rect 44272 43596 44324 43605
rect 19574 43494 19626 43546
rect 19638 43494 19690 43546
rect 19702 43494 19754 43546
rect 19766 43494 19818 43546
rect 19830 43494 19882 43546
rect 50294 43494 50346 43546
rect 50358 43494 50410 43546
rect 50422 43494 50474 43546
rect 50486 43494 50538 43546
rect 50550 43494 50602 43546
rect 40316 43435 40368 43444
rect 40316 43401 40331 43435
rect 40331 43401 40365 43435
rect 40365 43401 40368 43435
rect 40316 43392 40368 43401
rect 41236 43392 41288 43444
rect 41696 43435 41748 43444
rect 41696 43401 41705 43435
rect 41705 43401 41739 43435
rect 41739 43401 41748 43435
rect 41696 43392 41748 43401
rect 45560 43392 45612 43444
rect 45928 43392 45980 43444
rect 49424 43392 49476 43444
rect 53012 43392 53064 43444
rect 44180 43324 44232 43376
rect 47032 43324 47084 43376
rect 36452 43256 36504 43308
rect 38660 43256 38712 43308
rect 39488 43256 39540 43308
rect 37280 43231 37332 43240
rect 37280 43197 37289 43231
rect 37289 43197 37323 43231
rect 37323 43197 37332 43231
rect 37280 43188 37332 43197
rect 39856 43231 39908 43240
rect 39856 43197 39865 43231
rect 39865 43197 39899 43231
rect 39899 43197 39908 43231
rect 39856 43188 39908 43197
rect 45284 43299 45336 43308
rect 45284 43265 45293 43299
rect 45293 43265 45327 43299
rect 45327 43265 45336 43299
rect 45284 43256 45336 43265
rect 52460 43256 52512 43308
rect 52828 43256 52880 43308
rect 40500 43188 40552 43240
rect 45560 43231 45612 43240
rect 45560 43197 45569 43231
rect 45569 43197 45603 43231
rect 45603 43197 45612 43231
rect 45560 43188 45612 43197
rect 46940 43188 46992 43240
rect 49332 43231 49384 43240
rect 49332 43197 49341 43231
rect 49341 43197 49375 43231
rect 49375 43197 49384 43231
rect 49332 43188 49384 43197
rect 49700 43188 49752 43240
rect 50068 43231 50120 43240
rect 50068 43197 50077 43231
rect 50077 43197 50111 43231
rect 50111 43197 50120 43231
rect 50068 43188 50120 43197
rect 52920 43231 52972 43240
rect 52920 43197 52929 43231
rect 52929 43197 52963 43231
rect 52963 43197 52972 43231
rect 52920 43188 52972 43197
rect 4068 43052 4120 43104
rect 38660 43095 38712 43104
rect 38660 43061 38669 43095
rect 38669 43061 38703 43095
rect 38703 43061 38712 43095
rect 38660 43052 38712 43061
rect 41512 43052 41564 43104
rect 44180 43052 44232 43104
rect 45376 43052 45428 43104
rect 48136 43052 48188 43104
rect 53012 43120 53064 43172
rect 52736 43095 52788 43104
rect 52736 43061 52745 43095
rect 52745 43061 52779 43095
rect 52779 43061 52788 43095
rect 52736 43052 52788 43061
rect 4214 42950 4266 43002
rect 4278 42950 4330 43002
rect 4342 42950 4394 43002
rect 4406 42950 4458 43002
rect 4470 42950 4522 43002
rect 34934 42950 34986 43002
rect 34998 42950 35050 43002
rect 35062 42950 35114 43002
rect 35126 42950 35178 43002
rect 35190 42950 35242 43002
rect 38292 42848 38344 42900
rect 40500 42848 40552 42900
rect 45376 42891 45428 42900
rect 45376 42857 45385 42891
rect 45385 42857 45419 42891
rect 45419 42857 45428 42891
rect 45376 42848 45428 42857
rect 49332 42848 49384 42900
rect 38660 42712 38712 42764
rect 41512 42712 41564 42764
rect 45560 42712 45612 42764
rect 9588 42644 9640 42696
rect 36912 42687 36964 42696
rect 36912 42653 36946 42687
rect 36946 42653 36964 42687
rect 36912 42644 36964 42653
rect 37280 42576 37332 42628
rect 3976 42508 4028 42560
rect 41236 42508 41288 42560
rect 43076 42687 43128 42696
rect 43076 42653 43085 42687
rect 43085 42653 43119 42687
rect 43119 42653 43128 42687
rect 43076 42644 43128 42653
rect 47032 42780 47084 42832
rect 46020 42755 46072 42764
rect 46020 42721 46048 42755
rect 46048 42721 46072 42755
rect 48228 42755 48280 42764
rect 46020 42712 46072 42721
rect 48228 42721 48240 42755
rect 48240 42721 48274 42755
rect 48274 42721 48280 42755
rect 48228 42712 48280 42721
rect 45836 42687 45888 42696
rect 45836 42653 45845 42687
rect 45845 42653 45879 42687
rect 45879 42653 45888 42687
rect 45836 42644 45888 42653
rect 45928 42687 45980 42696
rect 45928 42653 45937 42687
rect 45937 42653 45971 42687
rect 45971 42653 45980 42687
rect 47768 42687 47820 42696
rect 45928 42644 45980 42653
rect 47768 42653 47777 42687
rect 47777 42653 47811 42687
rect 47811 42653 47820 42687
rect 47768 42644 47820 42653
rect 49424 42712 49476 42764
rect 48504 42687 48556 42696
rect 48504 42653 48513 42687
rect 48513 42653 48547 42687
rect 48547 42653 48556 42687
rect 48504 42644 48556 42653
rect 50068 42848 50120 42900
rect 50160 42712 50212 42764
rect 52644 42712 52696 42764
rect 43996 42576 44048 42628
rect 45560 42508 45612 42560
rect 46112 42619 46164 42628
rect 46112 42585 46121 42619
rect 46121 42585 46155 42619
rect 46155 42585 46164 42619
rect 46112 42576 46164 42585
rect 48136 42508 48188 42560
rect 52460 42644 52512 42696
rect 52552 42687 52604 42696
rect 52552 42653 52561 42687
rect 52561 42653 52595 42687
rect 52595 42653 52604 42687
rect 52552 42644 52604 42653
rect 56324 42644 56376 42696
rect 52092 42508 52144 42560
rect 57060 42576 57112 42628
rect 53656 42551 53708 42560
rect 53656 42517 53665 42551
rect 53665 42517 53699 42551
rect 53699 42517 53708 42551
rect 53656 42508 53708 42517
rect 19574 42406 19626 42458
rect 19638 42406 19690 42458
rect 19702 42406 19754 42458
rect 19766 42406 19818 42458
rect 19830 42406 19882 42458
rect 50294 42406 50346 42458
rect 50358 42406 50410 42458
rect 50422 42406 50474 42458
rect 50486 42406 50538 42458
rect 50550 42406 50602 42458
rect 44180 42347 44232 42356
rect 44180 42313 44189 42347
rect 44189 42313 44223 42347
rect 44223 42313 44232 42347
rect 44180 42304 44232 42313
rect 3976 42279 4028 42288
rect 3976 42245 3985 42279
rect 3985 42245 4019 42279
rect 4019 42245 4028 42279
rect 3976 42236 4028 42245
rect 45468 42304 45520 42356
rect 46112 42304 46164 42356
rect 47032 42304 47084 42356
rect 48504 42304 48556 42356
rect 45560 42236 45612 42288
rect 4160 42211 4212 42220
rect 4160 42177 4169 42211
rect 4169 42177 4203 42211
rect 4203 42177 4212 42211
rect 4160 42168 4212 42177
rect 44272 42211 44324 42220
rect 44272 42177 44281 42211
rect 44281 42177 44315 42211
rect 44315 42177 44324 42211
rect 44272 42168 44324 42177
rect 45100 42211 45152 42220
rect 45100 42177 45109 42211
rect 45109 42177 45143 42211
rect 45143 42177 45152 42211
rect 45100 42168 45152 42177
rect 2780 42143 2832 42152
rect 2780 42109 2789 42143
rect 2789 42109 2823 42143
rect 2823 42109 2832 42143
rect 2780 42100 2832 42109
rect 9588 42032 9640 42084
rect 33600 42032 33652 42084
rect 43996 42075 44048 42084
rect 43996 42041 44005 42075
rect 44005 42041 44039 42075
rect 44039 42041 44048 42075
rect 43996 42032 44048 42041
rect 49424 42304 49476 42356
rect 52000 42304 52052 42356
rect 52828 42304 52880 42356
rect 52920 42304 52972 42356
rect 53012 42211 53064 42220
rect 53012 42177 53021 42211
rect 53021 42177 53055 42211
rect 53055 42177 53064 42211
rect 53012 42168 53064 42177
rect 56876 42211 56928 42220
rect 56876 42177 56885 42211
rect 56885 42177 56919 42211
rect 56919 42177 56928 42211
rect 56876 42168 56928 42177
rect 49516 42143 49568 42152
rect 43076 41964 43128 42016
rect 49516 42109 49525 42143
rect 49525 42109 49559 42143
rect 49559 42109 49568 42143
rect 49516 42100 49568 42109
rect 49700 42100 49752 42152
rect 50068 42100 50120 42152
rect 50344 42100 50396 42152
rect 51080 42143 51132 42152
rect 51080 42109 51089 42143
rect 51089 42109 51123 42143
rect 51123 42109 51132 42143
rect 51080 42100 51132 42109
rect 51724 42100 51776 42152
rect 45744 41964 45796 42016
rect 47768 41964 47820 42016
rect 50068 41964 50120 42016
rect 56508 41964 56560 42016
rect 4214 41862 4266 41914
rect 4278 41862 4330 41914
rect 4342 41862 4394 41914
rect 4406 41862 4458 41914
rect 4470 41862 4522 41914
rect 34934 41862 34986 41914
rect 34998 41862 35050 41914
rect 35062 41862 35114 41914
rect 35126 41862 35178 41914
rect 35190 41862 35242 41914
rect 45100 41803 45152 41812
rect 45100 41769 45109 41803
rect 45109 41769 45143 41803
rect 45143 41769 45152 41803
rect 45100 41760 45152 41769
rect 46940 41760 46992 41812
rect 47124 41803 47176 41812
rect 47124 41769 47133 41803
rect 47133 41769 47167 41803
rect 47167 41769 47176 41803
rect 47124 41760 47176 41769
rect 52736 41803 52788 41812
rect 52736 41769 52745 41803
rect 52745 41769 52779 41803
rect 52779 41769 52788 41803
rect 52736 41760 52788 41769
rect 45744 41667 45796 41676
rect 45744 41633 45753 41667
rect 45753 41633 45787 41667
rect 45787 41633 45796 41667
rect 45744 41624 45796 41633
rect 51080 41624 51132 41676
rect 51724 41667 51776 41676
rect 51724 41633 51733 41667
rect 51733 41633 51767 41667
rect 51767 41633 51776 41667
rect 51724 41624 51776 41633
rect 56324 41667 56376 41676
rect 56324 41633 56333 41667
rect 56333 41633 56367 41667
rect 56367 41633 56376 41667
rect 56324 41624 56376 41633
rect 56508 41667 56560 41676
rect 56508 41633 56517 41667
rect 56517 41633 56551 41667
rect 56551 41633 56560 41667
rect 56508 41624 56560 41633
rect 58164 41667 58216 41676
rect 58164 41633 58173 41667
rect 58173 41633 58207 41667
rect 58207 41633 58216 41667
rect 58164 41624 58216 41633
rect 44180 41556 44232 41608
rect 46020 41599 46072 41608
rect 46020 41565 46054 41599
rect 46054 41565 46072 41599
rect 46020 41556 46072 41565
rect 47032 41488 47084 41540
rect 49516 41488 49568 41540
rect 53656 41556 53708 41608
rect 19574 41318 19626 41370
rect 19638 41318 19690 41370
rect 19702 41318 19754 41370
rect 19766 41318 19818 41370
rect 19830 41318 19882 41370
rect 50294 41318 50346 41370
rect 50358 41318 50410 41370
rect 50422 41318 50474 41370
rect 50486 41318 50538 41370
rect 50550 41318 50602 41370
rect 45836 41216 45888 41268
rect 45560 41123 45612 41132
rect 45560 41089 45569 41123
rect 45569 41089 45603 41123
rect 45603 41089 45612 41123
rect 45560 41080 45612 41089
rect 47124 41080 47176 41132
rect 4214 40774 4266 40826
rect 4278 40774 4330 40826
rect 4342 40774 4394 40826
rect 4406 40774 4458 40826
rect 4470 40774 4522 40826
rect 34934 40774 34986 40826
rect 34998 40774 35050 40826
rect 35062 40774 35114 40826
rect 35126 40774 35178 40826
rect 35190 40774 35242 40826
rect 19574 40230 19626 40282
rect 19638 40230 19690 40282
rect 19702 40230 19754 40282
rect 19766 40230 19818 40282
rect 19830 40230 19882 40282
rect 50294 40230 50346 40282
rect 50358 40230 50410 40282
rect 50422 40230 50474 40282
rect 50486 40230 50538 40282
rect 50550 40230 50602 40282
rect 4214 39686 4266 39738
rect 4278 39686 4330 39738
rect 4342 39686 4394 39738
rect 4406 39686 4458 39738
rect 4470 39686 4522 39738
rect 34934 39686 34986 39738
rect 34998 39686 35050 39738
rect 35062 39686 35114 39738
rect 35126 39686 35178 39738
rect 35190 39686 35242 39738
rect 19574 39142 19626 39194
rect 19638 39142 19690 39194
rect 19702 39142 19754 39194
rect 19766 39142 19818 39194
rect 19830 39142 19882 39194
rect 50294 39142 50346 39194
rect 50358 39142 50410 39194
rect 50422 39142 50474 39194
rect 50486 39142 50538 39194
rect 50550 39142 50602 39194
rect 4214 38598 4266 38650
rect 4278 38598 4330 38650
rect 4342 38598 4394 38650
rect 4406 38598 4458 38650
rect 4470 38598 4522 38650
rect 34934 38598 34986 38650
rect 34998 38598 35050 38650
rect 35062 38598 35114 38650
rect 35126 38598 35178 38650
rect 35190 38598 35242 38650
rect 19574 38054 19626 38106
rect 19638 38054 19690 38106
rect 19702 38054 19754 38106
rect 19766 38054 19818 38106
rect 19830 38054 19882 38106
rect 50294 38054 50346 38106
rect 50358 38054 50410 38106
rect 50422 38054 50474 38106
rect 50486 38054 50538 38106
rect 50550 38054 50602 38106
rect 4214 37510 4266 37562
rect 4278 37510 4330 37562
rect 4342 37510 4394 37562
rect 4406 37510 4458 37562
rect 4470 37510 4522 37562
rect 34934 37510 34986 37562
rect 34998 37510 35050 37562
rect 35062 37510 35114 37562
rect 35126 37510 35178 37562
rect 35190 37510 35242 37562
rect 19574 36966 19626 37018
rect 19638 36966 19690 37018
rect 19702 36966 19754 37018
rect 19766 36966 19818 37018
rect 19830 36966 19882 37018
rect 50294 36966 50346 37018
rect 50358 36966 50410 37018
rect 50422 36966 50474 37018
rect 50486 36966 50538 37018
rect 50550 36966 50602 37018
rect 4214 36422 4266 36474
rect 4278 36422 4330 36474
rect 4342 36422 4394 36474
rect 4406 36422 4458 36474
rect 4470 36422 4522 36474
rect 34934 36422 34986 36474
rect 34998 36422 35050 36474
rect 35062 36422 35114 36474
rect 35126 36422 35178 36474
rect 35190 36422 35242 36474
rect 19574 35878 19626 35930
rect 19638 35878 19690 35930
rect 19702 35878 19754 35930
rect 19766 35878 19818 35930
rect 19830 35878 19882 35930
rect 50294 35878 50346 35930
rect 50358 35878 50410 35930
rect 50422 35878 50474 35930
rect 50486 35878 50538 35930
rect 50550 35878 50602 35930
rect 4214 35334 4266 35386
rect 4278 35334 4330 35386
rect 4342 35334 4394 35386
rect 4406 35334 4458 35386
rect 4470 35334 4522 35386
rect 34934 35334 34986 35386
rect 34998 35334 35050 35386
rect 35062 35334 35114 35386
rect 35126 35334 35178 35386
rect 35190 35334 35242 35386
rect 2412 35071 2464 35080
rect 2412 35037 2421 35071
rect 2421 35037 2455 35071
rect 2455 35037 2464 35071
rect 2412 35028 2464 35037
rect 4620 35028 4672 35080
rect 9036 35028 9088 35080
rect 3792 34892 3844 34944
rect 19574 34790 19626 34842
rect 19638 34790 19690 34842
rect 19702 34790 19754 34842
rect 19766 34790 19818 34842
rect 19830 34790 19882 34842
rect 50294 34790 50346 34842
rect 50358 34790 50410 34842
rect 50422 34790 50474 34842
rect 50486 34790 50538 34842
rect 50550 34790 50602 34842
rect 2136 34663 2188 34672
rect 2136 34629 2145 34663
rect 2145 34629 2179 34663
rect 2179 34629 2188 34663
rect 2136 34620 2188 34629
rect 3792 34663 3844 34672
rect 3792 34629 3801 34663
rect 3801 34629 3835 34663
rect 3835 34629 3844 34663
rect 3792 34620 3844 34629
rect 2412 34484 2464 34536
rect 4214 34246 4266 34298
rect 4278 34246 4330 34298
rect 4342 34246 4394 34298
rect 4406 34246 4458 34298
rect 4470 34246 4522 34298
rect 34934 34246 34986 34298
rect 34998 34246 35050 34298
rect 35062 34246 35114 34298
rect 35126 34246 35178 34298
rect 35190 34246 35242 34298
rect 19574 33702 19626 33754
rect 19638 33702 19690 33754
rect 19702 33702 19754 33754
rect 19766 33702 19818 33754
rect 19830 33702 19882 33754
rect 50294 33702 50346 33754
rect 50358 33702 50410 33754
rect 50422 33702 50474 33754
rect 50486 33702 50538 33754
rect 50550 33702 50602 33754
rect 4214 33158 4266 33210
rect 4278 33158 4330 33210
rect 4342 33158 4394 33210
rect 4406 33158 4458 33210
rect 4470 33158 4522 33210
rect 34934 33158 34986 33210
rect 34998 33158 35050 33210
rect 35062 33158 35114 33210
rect 35126 33158 35178 33210
rect 35190 33158 35242 33210
rect 19574 32614 19626 32666
rect 19638 32614 19690 32666
rect 19702 32614 19754 32666
rect 19766 32614 19818 32666
rect 19830 32614 19882 32666
rect 50294 32614 50346 32666
rect 50358 32614 50410 32666
rect 50422 32614 50474 32666
rect 50486 32614 50538 32666
rect 50550 32614 50602 32666
rect 4214 32070 4266 32122
rect 4278 32070 4330 32122
rect 4342 32070 4394 32122
rect 4406 32070 4458 32122
rect 4470 32070 4522 32122
rect 34934 32070 34986 32122
rect 34998 32070 35050 32122
rect 35062 32070 35114 32122
rect 35126 32070 35178 32122
rect 35190 32070 35242 32122
rect 57060 31875 57112 31884
rect 57060 31841 57069 31875
rect 57069 31841 57103 31875
rect 57103 31841 57112 31875
rect 57060 31832 57112 31841
rect 58164 31807 58216 31816
rect 58164 31773 58173 31807
rect 58173 31773 58207 31807
rect 58207 31773 58216 31807
rect 58164 31764 58216 31773
rect 19574 31526 19626 31578
rect 19638 31526 19690 31578
rect 19702 31526 19754 31578
rect 19766 31526 19818 31578
rect 19830 31526 19882 31578
rect 50294 31526 50346 31578
rect 50358 31526 50410 31578
rect 50422 31526 50474 31578
rect 50486 31526 50538 31578
rect 50550 31526 50602 31578
rect 4214 30982 4266 31034
rect 4278 30982 4330 31034
rect 4342 30982 4394 31034
rect 4406 30982 4458 31034
rect 4470 30982 4522 31034
rect 34934 30982 34986 31034
rect 34998 30982 35050 31034
rect 35062 30982 35114 31034
rect 35126 30982 35178 31034
rect 35190 30982 35242 31034
rect 19574 30438 19626 30490
rect 19638 30438 19690 30490
rect 19702 30438 19754 30490
rect 19766 30438 19818 30490
rect 19830 30438 19882 30490
rect 50294 30438 50346 30490
rect 50358 30438 50410 30490
rect 50422 30438 50474 30490
rect 50486 30438 50538 30490
rect 50550 30438 50602 30490
rect 4214 29894 4266 29946
rect 4278 29894 4330 29946
rect 4342 29894 4394 29946
rect 4406 29894 4458 29946
rect 4470 29894 4522 29946
rect 34934 29894 34986 29946
rect 34998 29894 35050 29946
rect 35062 29894 35114 29946
rect 35126 29894 35178 29946
rect 35190 29894 35242 29946
rect 19574 29350 19626 29402
rect 19638 29350 19690 29402
rect 19702 29350 19754 29402
rect 19766 29350 19818 29402
rect 19830 29350 19882 29402
rect 50294 29350 50346 29402
rect 50358 29350 50410 29402
rect 50422 29350 50474 29402
rect 50486 29350 50538 29402
rect 50550 29350 50602 29402
rect 56968 29155 57020 29164
rect 56968 29121 56977 29155
rect 56977 29121 57011 29155
rect 57011 29121 57020 29155
rect 56968 29112 57020 29121
rect 57980 28976 58032 29028
rect 58164 28908 58216 28960
rect 4214 28806 4266 28858
rect 4278 28806 4330 28858
rect 4342 28806 4394 28858
rect 4406 28806 4458 28858
rect 4470 28806 4522 28858
rect 34934 28806 34986 28858
rect 34998 28806 35050 28858
rect 35062 28806 35114 28858
rect 35126 28806 35178 28858
rect 35190 28806 35242 28858
rect 57704 28611 57756 28620
rect 57704 28577 57713 28611
rect 57713 28577 57747 28611
rect 57747 28577 57756 28611
rect 57704 28568 57756 28577
rect 57980 28611 58032 28620
rect 57980 28577 57989 28611
rect 57989 28577 58023 28611
rect 58023 28577 58032 28611
rect 57980 28568 58032 28577
rect 58164 28611 58216 28620
rect 58164 28577 58173 28611
rect 58173 28577 58207 28611
rect 58207 28577 58216 28611
rect 58164 28568 58216 28577
rect 19574 28262 19626 28314
rect 19638 28262 19690 28314
rect 19702 28262 19754 28314
rect 19766 28262 19818 28314
rect 19830 28262 19882 28314
rect 50294 28262 50346 28314
rect 50358 28262 50410 28314
rect 50422 28262 50474 28314
rect 50486 28262 50538 28314
rect 50550 28262 50602 28314
rect 4214 27718 4266 27770
rect 4278 27718 4330 27770
rect 4342 27718 4394 27770
rect 4406 27718 4458 27770
rect 4470 27718 4522 27770
rect 34934 27718 34986 27770
rect 34998 27718 35050 27770
rect 35062 27718 35114 27770
rect 35126 27718 35178 27770
rect 35190 27718 35242 27770
rect 19574 27174 19626 27226
rect 19638 27174 19690 27226
rect 19702 27174 19754 27226
rect 19766 27174 19818 27226
rect 19830 27174 19882 27226
rect 50294 27174 50346 27226
rect 50358 27174 50410 27226
rect 50422 27174 50474 27226
rect 50486 27174 50538 27226
rect 50550 27174 50602 27226
rect 4214 26630 4266 26682
rect 4278 26630 4330 26682
rect 4342 26630 4394 26682
rect 4406 26630 4458 26682
rect 4470 26630 4522 26682
rect 34934 26630 34986 26682
rect 34998 26630 35050 26682
rect 35062 26630 35114 26682
rect 35126 26630 35178 26682
rect 35190 26630 35242 26682
rect 19574 26086 19626 26138
rect 19638 26086 19690 26138
rect 19702 26086 19754 26138
rect 19766 26086 19818 26138
rect 19830 26086 19882 26138
rect 50294 26086 50346 26138
rect 50358 26086 50410 26138
rect 50422 26086 50474 26138
rect 50486 26086 50538 26138
rect 50550 26086 50602 26138
rect 8208 26027 8260 26036
rect 8208 25993 8217 26027
rect 8217 25993 8251 26027
rect 8251 25993 8260 26027
rect 8208 25984 8260 25993
rect 8300 25891 8352 25900
rect 8300 25857 8309 25891
rect 8309 25857 8343 25891
rect 8343 25857 8352 25891
rect 8300 25848 8352 25857
rect 4214 25542 4266 25594
rect 4278 25542 4330 25594
rect 4342 25542 4394 25594
rect 4406 25542 4458 25594
rect 4470 25542 4522 25594
rect 34934 25542 34986 25594
rect 34998 25542 35050 25594
rect 35062 25542 35114 25594
rect 35126 25542 35178 25594
rect 35190 25542 35242 25594
rect 19574 24998 19626 25050
rect 19638 24998 19690 25050
rect 19702 24998 19754 25050
rect 19766 24998 19818 25050
rect 19830 24998 19882 25050
rect 50294 24998 50346 25050
rect 50358 24998 50410 25050
rect 50422 24998 50474 25050
rect 50486 24998 50538 25050
rect 50550 24998 50602 25050
rect 8300 24760 8352 24812
rect 57060 24803 57112 24812
rect 57060 24769 57069 24803
rect 57069 24769 57103 24803
rect 57103 24769 57112 24803
rect 57060 24760 57112 24769
rect 9588 24692 9640 24744
rect 56232 24735 56284 24744
rect 56232 24701 56241 24735
rect 56241 24701 56275 24735
rect 56275 24701 56284 24735
rect 56232 24692 56284 24701
rect 57796 24624 57848 24676
rect 56508 24556 56560 24608
rect 57888 24599 57940 24608
rect 57888 24565 57897 24599
rect 57897 24565 57931 24599
rect 57931 24565 57940 24599
rect 57888 24556 57940 24565
rect 4214 24454 4266 24506
rect 4278 24454 4330 24506
rect 4342 24454 4394 24506
rect 4406 24454 4458 24506
rect 4470 24454 4522 24506
rect 34934 24454 34986 24506
rect 34998 24454 35050 24506
rect 35062 24454 35114 24506
rect 35126 24454 35178 24506
rect 35190 24454 35242 24506
rect 57888 24284 57940 24336
rect 56508 24259 56560 24268
rect 56508 24225 56517 24259
rect 56517 24225 56551 24259
rect 56551 24225 56560 24259
rect 56508 24216 56560 24225
rect 58164 24259 58216 24268
rect 58164 24225 58173 24259
rect 58173 24225 58207 24259
rect 58207 24225 58216 24259
rect 58164 24216 58216 24225
rect 19574 23910 19626 23962
rect 19638 23910 19690 23962
rect 19702 23910 19754 23962
rect 19766 23910 19818 23962
rect 19830 23910 19882 23962
rect 50294 23910 50346 23962
rect 50358 23910 50410 23962
rect 50422 23910 50474 23962
rect 50486 23910 50538 23962
rect 50550 23910 50602 23962
rect 57060 23783 57112 23792
rect 57060 23749 57069 23783
rect 57069 23749 57103 23783
rect 57103 23749 57112 23783
rect 57060 23740 57112 23749
rect 55680 23468 55732 23520
rect 4214 23366 4266 23418
rect 4278 23366 4330 23418
rect 4342 23366 4394 23418
rect 4406 23366 4458 23418
rect 4470 23366 4522 23418
rect 34934 23366 34986 23418
rect 34998 23366 35050 23418
rect 35062 23366 35114 23418
rect 35126 23366 35178 23418
rect 35190 23366 35242 23418
rect 8300 23128 8352 23180
rect 7564 23060 7616 23112
rect 19574 22822 19626 22874
rect 19638 22822 19690 22874
rect 19702 22822 19754 22874
rect 19766 22822 19818 22874
rect 19830 22822 19882 22874
rect 50294 22822 50346 22874
rect 50358 22822 50410 22874
rect 50422 22822 50474 22874
rect 50486 22822 50538 22874
rect 50550 22822 50602 22874
rect 7564 22627 7616 22636
rect 7564 22593 7573 22627
rect 7573 22593 7607 22627
rect 7607 22593 7616 22627
rect 7564 22584 7616 22593
rect 8852 22423 8904 22432
rect 8852 22389 8861 22423
rect 8861 22389 8895 22423
rect 8895 22389 8904 22423
rect 8852 22380 8904 22389
rect 56968 22380 57020 22432
rect 4214 22278 4266 22330
rect 4278 22278 4330 22330
rect 4342 22278 4394 22330
rect 4406 22278 4458 22330
rect 4470 22278 4522 22330
rect 34934 22278 34986 22330
rect 34998 22278 35050 22330
rect 35062 22278 35114 22330
rect 35126 22278 35178 22330
rect 35190 22278 35242 22330
rect 19574 21734 19626 21786
rect 19638 21734 19690 21786
rect 19702 21734 19754 21786
rect 19766 21734 19818 21786
rect 19830 21734 19882 21786
rect 50294 21734 50346 21786
rect 50358 21734 50410 21786
rect 50422 21734 50474 21786
rect 50486 21734 50538 21786
rect 50550 21734 50602 21786
rect 4214 21190 4266 21242
rect 4278 21190 4330 21242
rect 4342 21190 4394 21242
rect 4406 21190 4458 21242
rect 4470 21190 4522 21242
rect 34934 21190 34986 21242
rect 34998 21190 35050 21242
rect 35062 21190 35114 21242
rect 35126 21190 35178 21242
rect 35190 21190 35242 21242
rect 19574 20646 19626 20698
rect 19638 20646 19690 20698
rect 19702 20646 19754 20698
rect 19766 20646 19818 20698
rect 19830 20646 19882 20698
rect 50294 20646 50346 20698
rect 50358 20646 50410 20698
rect 50422 20646 50474 20698
rect 50486 20646 50538 20698
rect 50550 20646 50602 20698
rect 4214 20102 4266 20154
rect 4278 20102 4330 20154
rect 4342 20102 4394 20154
rect 4406 20102 4458 20154
rect 4470 20102 4522 20154
rect 34934 20102 34986 20154
rect 34998 20102 35050 20154
rect 35062 20102 35114 20154
rect 35126 20102 35178 20154
rect 35190 20102 35242 20154
rect 19574 19558 19626 19610
rect 19638 19558 19690 19610
rect 19702 19558 19754 19610
rect 19766 19558 19818 19610
rect 19830 19558 19882 19610
rect 50294 19558 50346 19610
rect 50358 19558 50410 19610
rect 50422 19558 50474 19610
rect 50486 19558 50538 19610
rect 50550 19558 50602 19610
rect 56140 19320 56192 19372
rect 56508 19116 56560 19168
rect 57888 19159 57940 19168
rect 57888 19125 57897 19159
rect 57897 19125 57931 19159
rect 57931 19125 57940 19159
rect 57888 19116 57940 19125
rect 4214 19014 4266 19066
rect 4278 19014 4330 19066
rect 4342 19014 4394 19066
rect 4406 19014 4458 19066
rect 4470 19014 4522 19066
rect 34934 19014 34986 19066
rect 34998 19014 35050 19066
rect 35062 19014 35114 19066
rect 35126 19014 35178 19066
rect 35190 19014 35242 19066
rect 57888 18844 57940 18896
rect 56508 18819 56560 18828
rect 56508 18785 56517 18819
rect 56517 18785 56551 18819
rect 56551 18785 56560 18819
rect 56508 18776 56560 18785
rect 58164 18819 58216 18828
rect 58164 18785 58173 18819
rect 58173 18785 58207 18819
rect 58207 18785 58216 18819
rect 58164 18776 58216 18785
rect 19574 18470 19626 18522
rect 19638 18470 19690 18522
rect 19702 18470 19754 18522
rect 19766 18470 19818 18522
rect 19830 18470 19882 18522
rect 50294 18470 50346 18522
rect 50358 18470 50410 18522
rect 50422 18470 50474 18522
rect 50486 18470 50538 18522
rect 50550 18470 50602 18522
rect 4214 17926 4266 17978
rect 4278 17926 4330 17978
rect 4342 17926 4394 17978
rect 4406 17926 4458 17978
rect 4470 17926 4522 17978
rect 34934 17926 34986 17978
rect 34998 17926 35050 17978
rect 35062 17926 35114 17978
rect 35126 17926 35178 17978
rect 35190 17926 35242 17978
rect 19574 17382 19626 17434
rect 19638 17382 19690 17434
rect 19702 17382 19754 17434
rect 19766 17382 19818 17434
rect 19830 17382 19882 17434
rect 50294 17382 50346 17434
rect 50358 17382 50410 17434
rect 50422 17382 50474 17434
rect 50486 17382 50538 17434
rect 50550 17382 50602 17434
rect 4214 16838 4266 16890
rect 4278 16838 4330 16890
rect 4342 16838 4394 16890
rect 4406 16838 4458 16890
rect 4470 16838 4522 16890
rect 34934 16838 34986 16890
rect 34998 16838 35050 16890
rect 35062 16838 35114 16890
rect 35126 16838 35178 16890
rect 35190 16838 35242 16890
rect 19574 16294 19626 16346
rect 19638 16294 19690 16346
rect 19702 16294 19754 16346
rect 19766 16294 19818 16346
rect 19830 16294 19882 16346
rect 50294 16294 50346 16346
rect 50358 16294 50410 16346
rect 50422 16294 50474 16346
rect 50486 16294 50538 16346
rect 50550 16294 50602 16346
rect 4214 15750 4266 15802
rect 4278 15750 4330 15802
rect 4342 15750 4394 15802
rect 4406 15750 4458 15802
rect 4470 15750 4522 15802
rect 34934 15750 34986 15802
rect 34998 15750 35050 15802
rect 35062 15750 35114 15802
rect 35126 15750 35178 15802
rect 35190 15750 35242 15802
rect 19574 15206 19626 15258
rect 19638 15206 19690 15258
rect 19702 15206 19754 15258
rect 19766 15206 19818 15258
rect 19830 15206 19882 15258
rect 50294 15206 50346 15258
rect 50358 15206 50410 15258
rect 50422 15206 50474 15258
rect 50486 15206 50538 15258
rect 50550 15206 50602 15258
rect 4214 14662 4266 14714
rect 4278 14662 4330 14714
rect 4342 14662 4394 14714
rect 4406 14662 4458 14714
rect 4470 14662 4522 14714
rect 34934 14662 34986 14714
rect 34998 14662 35050 14714
rect 35062 14662 35114 14714
rect 35126 14662 35178 14714
rect 35190 14662 35242 14714
rect 19574 14118 19626 14170
rect 19638 14118 19690 14170
rect 19702 14118 19754 14170
rect 19766 14118 19818 14170
rect 19830 14118 19882 14170
rect 50294 14118 50346 14170
rect 50358 14118 50410 14170
rect 50422 14118 50474 14170
rect 50486 14118 50538 14170
rect 50550 14118 50602 14170
rect 4214 13574 4266 13626
rect 4278 13574 4330 13626
rect 4342 13574 4394 13626
rect 4406 13574 4458 13626
rect 4470 13574 4522 13626
rect 34934 13574 34986 13626
rect 34998 13574 35050 13626
rect 35062 13574 35114 13626
rect 35126 13574 35178 13626
rect 35190 13574 35242 13626
rect 19574 13030 19626 13082
rect 19638 13030 19690 13082
rect 19702 13030 19754 13082
rect 19766 13030 19818 13082
rect 19830 13030 19882 13082
rect 50294 13030 50346 13082
rect 50358 13030 50410 13082
rect 50422 13030 50474 13082
rect 50486 13030 50538 13082
rect 50550 13030 50602 13082
rect 4214 12486 4266 12538
rect 4278 12486 4330 12538
rect 4342 12486 4394 12538
rect 4406 12486 4458 12538
rect 4470 12486 4522 12538
rect 34934 12486 34986 12538
rect 34998 12486 35050 12538
rect 35062 12486 35114 12538
rect 35126 12486 35178 12538
rect 35190 12486 35242 12538
rect 56324 12180 56376 12232
rect 19574 11942 19626 11994
rect 19638 11942 19690 11994
rect 19702 11942 19754 11994
rect 19766 11942 19818 11994
rect 19830 11942 19882 11994
rect 50294 11942 50346 11994
rect 50358 11942 50410 11994
rect 50422 11942 50474 11994
rect 50486 11942 50538 11994
rect 50550 11942 50602 11994
rect 56968 11747 57020 11756
rect 56968 11713 56977 11747
rect 56977 11713 57011 11747
rect 57011 11713 57020 11747
rect 56968 11704 57020 11713
rect 56508 11500 56560 11552
rect 4214 11398 4266 11450
rect 4278 11398 4330 11450
rect 4342 11398 4394 11450
rect 4406 11398 4458 11450
rect 4470 11398 4522 11450
rect 34934 11398 34986 11450
rect 34998 11398 35050 11450
rect 35062 11398 35114 11450
rect 35126 11398 35178 11450
rect 35190 11398 35242 11450
rect 56324 11203 56376 11212
rect 56324 11169 56333 11203
rect 56333 11169 56367 11203
rect 56367 11169 56376 11203
rect 56324 11160 56376 11169
rect 56508 11203 56560 11212
rect 56508 11169 56517 11203
rect 56517 11169 56551 11203
rect 56551 11169 56560 11203
rect 56508 11160 56560 11169
rect 58164 11203 58216 11212
rect 58164 11169 58173 11203
rect 58173 11169 58207 11203
rect 58207 11169 58216 11203
rect 58164 11160 58216 11169
rect 8852 11092 8904 11144
rect 2136 10956 2188 11008
rect 19574 10854 19626 10906
rect 19638 10854 19690 10906
rect 19702 10854 19754 10906
rect 19766 10854 19818 10906
rect 19830 10854 19882 10906
rect 50294 10854 50346 10906
rect 50358 10854 50410 10906
rect 50422 10854 50474 10906
rect 50486 10854 50538 10906
rect 50550 10854 50602 10906
rect 2136 10727 2188 10736
rect 2136 10693 2145 10727
rect 2145 10693 2179 10727
rect 2179 10693 2188 10727
rect 2136 10684 2188 10693
rect 1952 10591 2004 10600
rect 1952 10557 1961 10591
rect 1961 10557 1995 10591
rect 1995 10557 2004 10591
rect 1952 10548 2004 10557
rect 2780 10591 2832 10600
rect 2780 10557 2789 10591
rect 2789 10557 2823 10591
rect 2823 10557 2832 10591
rect 2780 10548 2832 10557
rect 4214 10310 4266 10362
rect 4278 10310 4330 10362
rect 4342 10310 4394 10362
rect 4406 10310 4458 10362
rect 4470 10310 4522 10362
rect 34934 10310 34986 10362
rect 34998 10310 35050 10362
rect 35062 10310 35114 10362
rect 35126 10310 35178 10362
rect 35190 10310 35242 10362
rect 1952 10208 2004 10260
rect 19574 9766 19626 9818
rect 19638 9766 19690 9818
rect 19702 9766 19754 9818
rect 19766 9766 19818 9818
rect 19830 9766 19882 9818
rect 50294 9766 50346 9818
rect 50358 9766 50410 9818
rect 50422 9766 50474 9818
rect 50486 9766 50538 9818
rect 50550 9766 50602 9818
rect 4214 9222 4266 9274
rect 4278 9222 4330 9274
rect 4342 9222 4394 9274
rect 4406 9222 4458 9274
rect 4470 9222 4522 9274
rect 34934 9222 34986 9274
rect 34998 9222 35050 9274
rect 35062 9222 35114 9274
rect 35126 9222 35178 9274
rect 35190 9222 35242 9274
rect 57888 8984 57940 9036
rect 56508 8891 56560 8900
rect 56508 8857 56517 8891
rect 56517 8857 56551 8891
rect 56551 8857 56560 8891
rect 56508 8848 56560 8857
rect 58164 8891 58216 8900
rect 58164 8857 58173 8891
rect 58173 8857 58207 8891
rect 58207 8857 58216 8891
rect 58164 8848 58216 8857
rect 19574 8678 19626 8730
rect 19638 8678 19690 8730
rect 19702 8678 19754 8730
rect 19766 8678 19818 8730
rect 19830 8678 19882 8730
rect 50294 8678 50346 8730
rect 50358 8678 50410 8730
rect 50422 8678 50474 8730
rect 50486 8678 50538 8730
rect 50550 8678 50602 8730
rect 56508 8576 56560 8628
rect 56232 8440 56284 8492
rect 57888 8483 57940 8492
rect 57888 8449 57897 8483
rect 57897 8449 57931 8483
rect 57931 8449 57940 8483
rect 57888 8440 57940 8449
rect 4214 8134 4266 8186
rect 4278 8134 4330 8186
rect 4342 8134 4394 8186
rect 4406 8134 4458 8186
rect 4470 8134 4522 8186
rect 34934 8134 34986 8186
rect 34998 8134 35050 8186
rect 35062 8134 35114 8186
rect 35126 8134 35178 8186
rect 35190 8134 35242 8186
rect 19574 7590 19626 7642
rect 19638 7590 19690 7642
rect 19702 7590 19754 7642
rect 19766 7590 19818 7642
rect 19830 7590 19882 7642
rect 50294 7590 50346 7642
rect 50358 7590 50410 7642
rect 50422 7590 50474 7642
rect 50486 7590 50538 7642
rect 50550 7590 50602 7642
rect 4214 7046 4266 7098
rect 4278 7046 4330 7098
rect 4342 7046 4394 7098
rect 4406 7046 4458 7098
rect 4470 7046 4522 7098
rect 34934 7046 34986 7098
rect 34998 7046 35050 7098
rect 35062 7046 35114 7098
rect 35126 7046 35178 7098
rect 35190 7046 35242 7098
rect 19574 6502 19626 6554
rect 19638 6502 19690 6554
rect 19702 6502 19754 6554
rect 19766 6502 19818 6554
rect 19830 6502 19882 6554
rect 50294 6502 50346 6554
rect 50358 6502 50410 6554
rect 50422 6502 50474 6554
rect 50486 6502 50538 6554
rect 50550 6502 50602 6554
rect 4214 5958 4266 6010
rect 4278 5958 4330 6010
rect 4342 5958 4394 6010
rect 4406 5958 4458 6010
rect 4470 5958 4522 6010
rect 34934 5958 34986 6010
rect 34998 5958 35050 6010
rect 35062 5958 35114 6010
rect 35126 5958 35178 6010
rect 35190 5958 35242 6010
rect 19574 5414 19626 5466
rect 19638 5414 19690 5466
rect 19702 5414 19754 5466
rect 19766 5414 19818 5466
rect 19830 5414 19882 5466
rect 50294 5414 50346 5466
rect 50358 5414 50410 5466
rect 50422 5414 50474 5466
rect 50486 5414 50538 5466
rect 50550 5414 50602 5466
rect 1952 4972 2004 5024
rect 4214 4870 4266 4922
rect 4278 4870 4330 4922
rect 4342 4870 4394 4922
rect 4406 4870 4458 4922
rect 4470 4870 4522 4922
rect 34934 4870 34986 4922
rect 34998 4870 35050 4922
rect 35062 4870 35114 4922
rect 35126 4870 35178 4922
rect 35190 4870 35242 4922
rect 2504 4607 2556 4616
rect 2504 4573 2513 4607
rect 2513 4573 2547 4607
rect 2547 4573 2556 4607
rect 2504 4564 2556 4573
rect 8208 4564 8260 4616
rect 56324 4607 56376 4616
rect 56324 4573 56333 4607
rect 56333 4573 56367 4607
rect 56367 4573 56376 4607
rect 56324 4564 56376 4573
rect 56508 4539 56560 4548
rect 56508 4505 56517 4539
rect 56517 4505 56551 4539
rect 56551 4505 56560 4539
rect 56508 4496 56560 4505
rect 59268 4496 59320 4548
rect 2136 4428 2188 4480
rect 19574 4326 19626 4378
rect 19638 4326 19690 4378
rect 19702 4326 19754 4378
rect 19766 4326 19818 4378
rect 19830 4326 19882 4378
rect 50294 4326 50346 4378
rect 50358 4326 50410 4378
rect 50422 4326 50474 4378
rect 50486 4326 50538 4378
rect 50550 4326 50602 4378
rect 2136 4199 2188 4208
rect 2136 4165 2145 4199
rect 2145 4165 2179 4199
rect 2179 4165 2188 4199
rect 2136 4156 2188 4165
rect 1952 4131 2004 4140
rect 1952 4097 1961 4131
rect 1961 4097 1995 4131
rect 1995 4097 2004 4131
rect 1952 4088 2004 4097
rect 7564 4131 7616 4140
rect 7564 4097 7573 4131
rect 7573 4097 7607 4131
rect 7607 4097 7616 4131
rect 7564 4088 7616 4097
rect 57796 4088 57848 4140
rect 2780 4063 2832 4072
rect 2780 4029 2789 4063
rect 2789 4029 2823 4063
rect 2823 4029 2832 4063
rect 2780 4020 2832 4029
rect 4712 4020 4764 4072
rect 51448 4020 51500 4072
rect 57336 4063 57388 4072
rect 4068 3884 4120 3936
rect 20628 3884 20680 3936
rect 51540 3927 51592 3936
rect 51540 3893 51549 3927
rect 51549 3893 51583 3927
rect 51583 3893 51592 3927
rect 51540 3884 51592 3893
rect 54484 3927 54536 3936
rect 54484 3893 54493 3927
rect 54493 3893 54527 3927
rect 54527 3893 54536 3927
rect 54484 3884 54536 3893
rect 57336 4029 57345 4063
rect 57345 4029 57379 4063
rect 57379 4029 57388 4063
rect 57336 4020 57388 4029
rect 57244 3884 57296 3936
rect 4214 3782 4266 3834
rect 4278 3782 4330 3834
rect 4342 3782 4394 3834
rect 4406 3782 4458 3834
rect 4470 3782 4522 3834
rect 34934 3782 34986 3834
rect 34998 3782 35050 3834
rect 35062 3782 35114 3834
rect 35126 3782 35178 3834
rect 35190 3782 35242 3834
rect 56508 3680 56560 3732
rect 4068 3587 4120 3596
rect 4068 3553 4077 3587
rect 4077 3553 4111 3587
rect 4111 3553 4120 3587
rect 4068 3544 4120 3553
rect 4620 3587 4672 3596
rect 4620 3553 4629 3587
rect 4629 3553 4663 3587
rect 4663 3553 4672 3587
rect 4620 3544 4672 3553
rect 14188 3544 14240 3596
rect 7564 3519 7616 3528
rect 7564 3485 7573 3519
rect 7573 3485 7607 3519
rect 7607 3485 7616 3519
rect 7564 3476 7616 3485
rect 14464 3519 14516 3528
rect 14464 3485 14473 3519
rect 14473 3485 14507 3519
rect 14507 3485 14516 3519
rect 14464 3476 14516 3485
rect 4252 3451 4304 3460
rect 4252 3417 4261 3451
rect 4261 3417 4295 3451
rect 4295 3417 4304 3451
rect 4252 3408 4304 3417
rect 8208 3451 8260 3460
rect 8208 3417 8217 3451
rect 8217 3417 8251 3451
rect 8251 3417 8260 3451
rect 8208 3408 8260 3417
rect 15476 3408 15528 3460
rect 18696 3519 18748 3528
rect 18696 3485 18705 3519
rect 18705 3485 18739 3519
rect 18739 3485 18748 3519
rect 20628 3519 20680 3528
rect 18696 3476 18748 3485
rect 20628 3485 20637 3519
rect 20637 3485 20671 3519
rect 20671 3485 20680 3519
rect 20628 3476 20680 3485
rect 56784 3612 56836 3664
rect 45192 3544 45244 3596
rect 51540 3587 51592 3596
rect 51540 3553 51549 3587
rect 51549 3553 51583 3587
rect 51583 3553 51592 3587
rect 51540 3544 51592 3553
rect 52184 3587 52236 3596
rect 52184 3553 52193 3587
rect 52193 3553 52227 3587
rect 52227 3553 52236 3587
rect 52184 3544 52236 3553
rect 57888 3587 57940 3596
rect 57888 3553 57897 3587
rect 57897 3553 57931 3587
rect 57931 3553 57940 3587
rect 57888 3544 57940 3553
rect 44640 3476 44692 3528
rect 16764 3408 16816 3460
rect 18420 3408 18472 3460
rect 20812 3451 20864 3460
rect 20812 3417 20821 3451
rect 20821 3417 20855 3451
rect 20855 3417 20864 3451
rect 20812 3408 20864 3417
rect 21272 3408 21324 3460
rect 51724 3451 51776 3460
rect 51724 3417 51733 3451
rect 51733 3417 51767 3451
rect 51767 3417 51776 3451
rect 51724 3408 51776 3417
rect 50160 3340 50212 3392
rect 55680 3519 55732 3528
rect 55680 3485 55689 3519
rect 55689 3485 55723 3519
rect 55723 3485 55732 3519
rect 55680 3476 55732 3485
rect 56324 3519 56376 3528
rect 56324 3485 56333 3519
rect 56333 3485 56367 3519
rect 56367 3485 56376 3519
rect 56324 3476 56376 3485
rect 56876 3408 56928 3460
rect 54668 3383 54720 3392
rect 54668 3349 54677 3383
rect 54677 3349 54711 3383
rect 54711 3349 54720 3383
rect 54668 3340 54720 3349
rect 19574 3238 19626 3290
rect 19638 3238 19690 3290
rect 19702 3238 19754 3290
rect 19766 3238 19818 3290
rect 19830 3238 19882 3290
rect 50294 3238 50346 3290
rect 50358 3238 50410 3290
rect 50422 3238 50474 3290
rect 50486 3238 50538 3290
rect 50550 3238 50602 3290
rect 4252 3179 4304 3188
rect 4252 3145 4261 3179
rect 4261 3145 4295 3179
rect 4295 3145 4304 3179
rect 4252 3136 4304 3145
rect 15476 3179 15528 3188
rect 15476 3145 15485 3179
rect 15485 3145 15519 3179
rect 15519 3145 15528 3179
rect 15476 3136 15528 3145
rect 18420 3179 18472 3188
rect 18420 3145 18429 3179
rect 18429 3145 18463 3179
rect 18463 3145 18472 3179
rect 18420 3136 18472 3145
rect 20812 3179 20864 3188
rect 20812 3145 20821 3179
rect 20821 3145 20855 3179
rect 20855 3145 20864 3179
rect 20812 3136 20864 3145
rect 51724 3136 51776 3188
rect 4712 3000 4764 3052
rect 14464 3043 14516 3052
rect 14464 3009 14473 3043
rect 14473 3009 14507 3043
rect 14507 3009 14516 3043
rect 14464 3000 14516 3009
rect 18696 3068 18748 3120
rect 56140 3136 56192 3188
rect 56876 3179 56928 3188
rect 56876 3145 56885 3179
rect 56885 3145 56919 3179
rect 56919 3145 56928 3179
rect 56876 3136 56928 3145
rect 54668 3111 54720 3120
rect 44640 3043 44692 3052
rect 44640 3009 44649 3043
rect 44649 3009 44683 3043
rect 44683 3009 44692 3043
rect 44640 3000 44692 3009
rect 50160 2864 50212 2916
rect 51448 3000 51500 3052
rect 54668 3077 54677 3111
rect 54677 3077 54711 3111
rect 54711 3077 54720 3111
rect 54668 3068 54720 3077
rect 56324 3068 56376 3120
rect 54484 3043 54536 3052
rect 54484 3009 54493 3043
rect 54493 3009 54527 3043
rect 54527 3009 54536 3043
rect 54484 3000 54536 3009
rect 56784 3043 56836 3052
rect 56784 3009 56793 3043
rect 56793 3009 56827 3043
rect 56827 3009 56836 3043
rect 56784 3000 56836 3009
rect 54760 2932 54812 2984
rect 56232 2864 56284 2916
rect 4214 2694 4266 2746
rect 4278 2694 4330 2746
rect 4342 2694 4394 2746
rect 4406 2694 4458 2746
rect 4470 2694 4522 2746
rect 34934 2694 34986 2746
rect 34998 2694 35050 2746
rect 35062 2694 35114 2746
rect 35126 2694 35178 2746
rect 35190 2694 35242 2746
rect 7564 2635 7616 2644
rect 7564 2601 7573 2635
rect 7573 2601 7607 2635
rect 7607 2601 7616 2635
rect 7564 2592 7616 2601
rect 57336 2592 57388 2644
rect 56416 2524 56468 2576
rect 23848 2388 23900 2440
rect 7104 2320 7156 2372
rect 41512 2320 41564 2372
rect 19574 2150 19626 2202
rect 19638 2150 19690 2202
rect 19702 2150 19754 2202
rect 19766 2150 19818 2202
rect 19830 2150 19882 2202
rect 50294 2150 50346 2202
rect 50358 2150 50410 2202
rect 50422 2150 50474 2202
rect 50486 2150 50538 2202
rect 50550 2150 50602 2202
<< metal2 >>
rect 634 59200 746 60000
rect 2566 59200 2678 60000
rect 5142 59200 5254 60000
rect 7718 59200 7830 60000
rect 9650 59200 9762 60000
rect 12226 59200 12338 60000
rect 14802 59200 14914 60000
rect 17378 59200 17490 60000
rect 19310 59200 19422 60000
rect 21886 59200 21998 60000
rect 24462 59200 24574 60000
rect 26394 59200 26506 60000
rect 28970 59200 29082 60000
rect 31546 59200 31658 60000
rect 34122 59200 34234 60000
rect 36054 59200 36166 60000
rect 38630 59200 38742 60000
rect 41206 59200 41318 60000
rect 43138 59200 43250 60000
rect 45714 59200 45826 60000
rect 48290 59200 48402 60000
rect 50866 59200 50978 60000
rect 52798 59200 52910 60000
rect 55374 59200 55486 60000
rect 57950 59200 58062 60000
rect 59882 59200 59994 60000
rect 676 56438 704 59200
rect 4214 57148 4522 57168
rect 4214 57146 4220 57148
rect 4276 57146 4300 57148
rect 4356 57146 4380 57148
rect 4436 57146 4460 57148
rect 4516 57146 4522 57148
rect 4276 57094 4278 57146
rect 4458 57094 4460 57146
rect 4214 57092 4220 57094
rect 4276 57092 4300 57094
rect 4356 57092 4380 57094
rect 4436 57092 4460 57094
rect 4516 57092 4522 57094
rect 4214 57072 4522 57092
rect 664 56432 716 56438
rect 664 56374 716 56380
rect 7760 56302 7788 59200
rect 8484 56840 8536 56846
rect 8484 56782 8536 56788
rect 8944 56840 8996 56846
rect 8944 56782 8996 56788
rect 8496 56370 8524 56782
rect 8956 56370 8984 56782
rect 8484 56364 8536 56370
rect 8484 56306 8536 56312
rect 8944 56364 8996 56370
rect 8944 56306 8996 56312
rect 9692 56302 9720 59200
rect 19574 57692 19882 57712
rect 19574 57690 19580 57692
rect 19636 57690 19660 57692
rect 19716 57690 19740 57692
rect 19796 57690 19820 57692
rect 19876 57690 19882 57692
rect 19636 57638 19638 57690
rect 19818 57638 19820 57690
rect 19574 57636 19580 57638
rect 19636 57636 19660 57638
rect 19716 57636 19740 57638
rect 19796 57636 19820 57638
rect 19876 57636 19882 57638
rect 19574 57616 19882 57636
rect 25964 56840 26016 56846
rect 25964 56782 26016 56788
rect 19574 56604 19882 56624
rect 19574 56602 19580 56604
rect 19636 56602 19660 56604
rect 19716 56602 19740 56604
rect 19796 56602 19820 56604
rect 19876 56602 19882 56604
rect 19636 56550 19638 56602
rect 19818 56550 19820 56602
rect 19574 56548 19580 56550
rect 19636 56548 19660 56550
rect 19716 56548 19740 56550
rect 19796 56548 19820 56550
rect 19876 56548 19882 56550
rect 19574 56528 19882 56548
rect 7748 56296 7800 56302
rect 7748 56238 7800 56244
rect 8208 56296 8260 56302
rect 8208 56238 8260 56244
rect 9128 56296 9180 56302
rect 9128 56238 9180 56244
rect 9680 56296 9732 56302
rect 9680 56238 9732 56244
rect 4214 56060 4522 56080
rect 4214 56058 4220 56060
rect 4276 56058 4300 56060
rect 4356 56058 4380 56060
rect 4436 56058 4460 56060
rect 4516 56058 4522 56060
rect 4276 56006 4278 56058
rect 4458 56006 4460 56058
rect 4214 56004 4220 56006
rect 4276 56004 4300 56006
rect 4356 56004 4380 56006
rect 4436 56004 4460 56006
rect 4516 56004 4522 56006
rect 4214 55984 4522 56004
rect 2778 55176 2834 55185
rect 2778 55111 2834 55120
rect 1952 54664 2004 54670
rect 1952 54606 2004 54612
rect 1964 54194 1992 54606
rect 1952 54188 2004 54194
rect 1952 54130 2004 54136
rect 2792 54126 2820 55111
rect 4214 54972 4522 54992
rect 4214 54970 4220 54972
rect 4276 54970 4300 54972
rect 4356 54970 4380 54972
rect 4436 54970 4460 54972
rect 4516 54970 4522 54972
rect 4276 54918 4278 54970
rect 4458 54918 4460 54970
rect 4214 54916 4220 54918
rect 4276 54916 4300 54918
rect 4356 54916 4380 54918
rect 4436 54916 4460 54918
rect 4516 54916 4522 54918
rect 4214 54896 4522 54916
rect 2136 54120 2188 54126
rect 2136 54062 2188 54068
rect 2780 54120 2832 54126
rect 2780 54062 2832 54068
rect 2148 53786 2176 54062
rect 4214 53884 4522 53904
rect 4214 53882 4220 53884
rect 4276 53882 4300 53884
rect 4356 53882 4380 53884
rect 4436 53882 4460 53884
rect 4516 53882 4522 53884
rect 4276 53830 4278 53882
rect 4458 53830 4460 53882
rect 4214 53828 4220 53830
rect 4276 53828 4300 53830
rect 4356 53828 4380 53830
rect 4436 53828 4460 53830
rect 4516 53828 4522 53830
rect 4214 53808 4522 53828
rect 2136 53780 2188 53786
rect 2136 53722 2188 53728
rect 2596 53576 2648 53582
rect 2596 53518 2648 53524
rect 1952 49768 2004 49774
rect 1952 49710 2004 49716
rect 2136 49768 2188 49774
rect 2136 49710 2188 49716
rect 1964 49434 1992 49710
rect 1952 49428 2004 49434
rect 1952 49370 2004 49376
rect 2148 48890 2176 49710
rect 2136 48884 2188 48890
rect 2136 48826 2188 48832
rect 2504 48748 2556 48754
rect 2504 48690 2556 48696
rect 1952 48136 2004 48142
rect 1952 48078 2004 48084
rect 1964 47666 1992 48078
rect 1952 47660 2004 47666
rect 1952 47602 2004 47608
rect 2412 47592 2464 47598
rect 2412 47534 2464 47540
rect 2424 47258 2452 47534
rect 2412 47252 2464 47258
rect 2412 47194 2464 47200
rect 1952 45280 2004 45286
rect 1952 45222 2004 45228
rect 1964 44402 1992 45222
rect 2516 44878 2544 48690
rect 2608 47054 2636 53518
rect 4214 52796 4522 52816
rect 4214 52794 4220 52796
rect 4276 52794 4300 52796
rect 4356 52794 4380 52796
rect 4436 52794 4460 52796
rect 4516 52794 4522 52796
rect 4276 52742 4278 52794
rect 4458 52742 4460 52794
rect 4214 52740 4220 52742
rect 4276 52740 4300 52742
rect 4356 52740 4380 52742
rect 4436 52740 4460 52742
rect 4516 52740 4522 52742
rect 4214 52720 4522 52740
rect 4214 51708 4522 51728
rect 4214 51706 4220 51708
rect 4276 51706 4300 51708
rect 4356 51706 4380 51708
rect 4436 51706 4460 51708
rect 4516 51706 4522 51708
rect 4276 51654 4278 51706
rect 4458 51654 4460 51706
rect 4214 51652 4220 51654
rect 4276 51652 4300 51654
rect 4356 51652 4380 51654
rect 4436 51652 4460 51654
rect 4516 51652 4522 51654
rect 4214 51632 4522 51652
rect 4214 50620 4522 50640
rect 4214 50618 4220 50620
rect 4276 50618 4300 50620
rect 4356 50618 4380 50620
rect 4436 50618 4460 50620
rect 4516 50618 4522 50620
rect 4276 50566 4278 50618
rect 4458 50566 4460 50618
rect 4214 50564 4220 50566
rect 4276 50564 4300 50566
rect 4356 50564 4380 50566
rect 4436 50564 4460 50566
rect 4516 50564 4522 50566
rect 4214 50544 4522 50564
rect 2778 50416 2834 50425
rect 2778 50351 2834 50360
rect 2792 49774 2820 50351
rect 2780 49768 2832 49774
rect 2780 49710 2832 49716
rect 4214 49532 4522 49552
rect 4214 49530 4220 49532
rect 4276 49530 4300 49532
rect 4356 49530 4380 49532
rect 4436 49530 4460 49532
rect 4516 49530 4522 49532
rect 4276 49478 4278 49530
rect 4458 49478 4460 49530
rect 4214 49476 4220 49478
rect 4276 49476 4300 49478
rect 4356 49476 4380 49478
rect 4436 49476 4460 49478
rect 4516 49476 4522 49478
rect 4214 49456 4522 49476
rect 4214 48444 4522 48464
rect 4214 48442 4220 48444
rect 4276 48442 4300 48444
rect 4356 48442 4380 48444
rect 4436 48442 4460 48444
rect 4516 48442 4522 48444
rect 4276 48390 4278 48442
rect 4458 48390 4460 48442
rect 4214 48388 4220 48390
rect 4276 48388 4300 48390
rect 4356 48388 4380 48390
rect 4436 48388 4460 48390
rect 4516 48388 4522 48390
rect 4214 48368 4522 48388
rect 2778 47696 2834 47705
rect 2778 47631 2834 47640
rect 2792 47598 2820 47631
rect 2780 47592 2832 47598
rect 2780 47534 2832 47540
rect 4214 47356 4522 47376
rect 4214 47354 4220 47356
rect 4276 47354 4300 47356
rect 4356 47354 4380 47356
rect 4436 47354 4460 47356
rect 4516 47354 4522 47356
rect 4276 47302 4278 47354
rect 4458 47302 4460 47354
rect 4214 47300 4220 47302
rect 4276 47300 4300 47302
rect 4356 47300 4380 47302
rect 4436 47300 4460 47302
rect 4516 47300 4522 47302
rect 4214 47280 4522 47300
rect 2596 47048 2648 47054
rect 2596 46990 2648 46996
rect 4214 46268 4522 46288
rect 4214 46266 4220 46268
rect 4276 46266 4300 46268
rect 4356 46266 4380 46268
rect 4436 46266 4460 46268
rect 4516 46266 4522 46268
rect 4276 46214 4278 46266
rect 4458 46214 4460 46266
rect 4214 46212 4220 46214
rect 4276 46212 4300 46214
rect 4356 46212 4380 46214
rect 4436 46212 4460 46214
rect 4516 46212 4522 46214
rect 4214 46192 4522 46212
rect 4214 45180 4522 45200
rect 4214 45178 4220 45180
rect 4276 45178 4300 45180
rect 4356 45178 4380 45180
rect 4436 45178 4460 45180
rect 4516 45178 4522 45180
rect 4276 45126 4278 45178
rect 4458 45126 4460 45178
rect 4214 45124 4220 45126
rect 4276 45124 4300 45126
rect 4356 45124 4380 45126
rect 4436 45124 4460 45126
rect 4516 45124 4522 45126
rect 4214 45104 4522 45124
rect 2778 44976 2834 44985
rect 2778 44911 2834 44920
rect 2504 44872 2556 44878
rect 2504 44814 2556 44820
rect 2136 44736 2188 44742
rect 2136 44678 2188 44684
rect 2148 44470 2176 44678
rect 2136 44464 2188 44470
rect 2136 44406 2188 44412
rect 1952 44396 2004 44402
rect 1952 44338 2004 44344
rect 2412 35080 2464 35086
rect 2412 35022 2464 35028
rect 2134 34776 2190 34785
rect 2134 34711 2190 34720
rect 2148 34678 2176 34711
rect 2136 34672 2188 34678
rect 2136 34614 2188 34620
rect 2424 34542 2452 35022
rect 2412 34536 2464 34542
rect 2412 34478 2464 34484
rect 2136 11008 2188 11014
rect 2136 10950 2188 10956
rect 2148 10742 2176 10950
rect 2136 10736 2188 10742
rect 2136 10678 2188 10684
rect 1952 10600 2004 10606
rect 1952 10542 2004 10548
rect 1964 10266 1992 10542
rect 1952 10260 2004 10266
rect 1952 10202 2004 10208
rect 1952 5024 2004 5030
rect 1952 4966 2004 4972
rect 1964 4146 1992 4966
rect 2516 4622 2544 44814
rect 2792 44334 2820 44911
rect 2780 44328 2832 44334
rect 2780 44270 2832 44276
rect 4214 44092 4522 44112
rect 4214 44090 4220 44092
rect 4276 44090 4300 44092
rect 4356 44090 4380 44092
rect 4436 44090 4460 44092
rect 4516 44090 4522 44092
rect 4276 44038 4278 44090
rect 4458 44038 4460 44090
rect 4214 44036 4220 44038
rect 4276 44036 4300 44038
rect 4356 44036 4380 44038
rect 4436 44036 4460 44038
rect 4516 44036 4522 44038
rect 4214 44016 4522 44036
rect 4068 43104 4120 43110
rect 4068 43046 4120 43052
rect 2778 42936 2834 42945
rect 2778 42871 2834 42880
rect 2792 42158 2820 42871
rect 4080 42786 4108 43046
rect 4214 43004 4522 43024
rect 4214 43002 4220 43004
rect 4276 43002 4300 43004
rect 4356 43002 4380 43004
rect 4436 43002 4460 43004
rect 4516 43002 4522 43004
rect 4276 42950 4278 43002
rect 4458 42950 4460 43002
rect 4214 42948 4220 42950
rect 4276 42948 4300 42950
rect 4356 42948 4380 42950
rect 4436 42948 4460 42950
rect 4516 42948 4522 42950
rect 4214 42928 4522 42948
rect 4080 42758 4200 42786
rect 3976 42560 4028 42566
rect 3976 42502 4028 42508
rect 3988 42294 4016 42502
rect 3976 42288 4028 42294
rect 3976 42230 4028 42236
rect 4172 42226 4200 42758
rect 4160 42220 4212 42226
rect 4160 42162 4212 42168
rect 2780 42152 2832 42158
rect 2780 42094 2832 42100
rect 4214 41916 4522 41936
rect 4214 41914 4220 41916
rect 4276 41914 4300 41916
rect 4356 41914 4380 41916
rect 4436 41914 4460 41916
rect 4516 41914 4522 41916
rect 4276 41862 4278 41914
rect 4458 41862 4460 41914
rect 4214 41860 4220 41862
rect 4276 41860 4300 41862
rect 4356 41860 4380 41862
rect 4436 41860 4460 41862
rect 4516 41860 4522 41862
rect 4214 41840 4522 41860
rect 4214 40828 4522 40848
rect 4214 40826 4220 40828
rect 4276 40826 4300 40828
rect 4356 40826 4380 40828
rect 4436 40826 4460 40828
rect 4516 40826 4522 40828
rect 4276 40774 4278 40826
rect 4458 40774 4460 40826
rect 4214 40772 4220 40774
rect 4276 40772 4300 40774
rect 4356 40772 4380 40774
rect 4436 40772 4460 40774
rect 4516 40772 4522 40774
rect 4214 40752 4522 40772
rect 4214 39740 4522 39760
rect 4214 39738 4220 39740
rect 4276 39738 4300 39740
rect 4356 39738 4380 39740
rect 4436 39738 4460 39740
rect 4516 39738 4522 39740
rect 4276 39686 4278 39738
rect 4458 39686 4460 39738
rect 4214 39684 4220 39686
rect 4276 39684 4300 39686
rect 4356 39684 4380 39686
rect 4436 39684 4460 39686
rect 4516 39684 4522 39686
rect 4214 39664 4522 39684
rect 4214 38652 4522 38672
rect 4214 38650 4220 38652
rect 4276 38650 4300 38652
rect 4356 38650 4380 38652
rect 4436 38650 4460 38652
rect 4516 38650 4522 38652
rect 4276 38598 4278 38650
rect 4458 38598 4460 38650
rect 4214 38596 4220 38598
rect 4276 38596 4300 38598
rect 4356 38596 4380 38598
rect 4436 38596 4460 38598
rect 4516 38596 4522 38598
rect 4214 38576 4522 38596
rect 4214 37564 4522 37584
rect 4214 37562 4220 37564
rect 4276 37562 4300 37564
rect 4356 37562 4380 37564
rect 4436 37562 4460 37564
rect 4516 37562 4522 37564
rect 4276 37510 4278 37562
rect 4458 37510 4460 37562
rect 4214 37508 4220 37510
rect 4276 37508 4300 37510
rect 4356 37508 4380 37510
rect 4436 37508 4460 37510
rect 4516 37508 4522 37510
rect 4214 37488 4522 37508
rect 4214 36476 4522 36496
rect 4214 36474 4220 36476
rect 4276 36474 4300 36476
rect 4356 36474 4380 36476
rect 4436 36474 4460 36476
rect 4516 36474 4522 36476
rect 4276 36422 4278 36474
rect 4458 36422 4460 36474
rect 4214 36420 4220 36422
rect 4276 36420 4300 36422
rect 4356 36420 4380 36422
rect 4436 36420 4460 36422
rect 4516 36420 4522 36422
rect 4214 36400 4522 36420
rect 4214 35388 4522 35408
rect 4214 35386 4220 35388
rect 4276 35386 4300 35388
rect 4356 35386 4380 35388
rect 4436 35386 4460 35388
rect 4516 35386 4522 35388
rect 4276 35334 4278 35386
rect 4458 35334 4460 35386
rect 4214 35332 4220 35334
rect 4276 35332 4300 35334
rect 4356 35332 4380 35334
rect 4436 35332 4460 35334
rect 4516 35332 4522 35334
rect 4214 35312 4522 35332
rect 4620 35080 4672 35086
rect 4620 35022 4672 35028
rect 3792 34944 3844 34950
rect 3792 34886 3844 34892
rect 3804 34678 3832 34886
rect 3792 34672 3844 34678
rect 3792 34614 3844 34620
rect 4214 34300 4522 34320
rect 4214 34298 4220 34300
rect 4276 34298 4300 34300
rect 4356 34298 4380 34300
rect 4436 34298 4460 34300
rect 4516 34298 4522 34300
rect 4276 34246 4278 34298
rect 4458 34246 4460 34298
rect 4214 34244 4220 34246
rect 4276 34244 4300 34246
rect 4356 34244 4380 34246
rect 4436 34244 4460 34246
rect 4516 34244 4522 34246
rect 4214 34224 4522 34244
rect 4214 33212 4522 33232
rect 4214 33210 4220 33212
rect 4276 33210 4300 33212
rect 4356 33210 4380 33212
rect 4436 33210 4460 33212
rect 4516 33210 4522 33212
rect 4276 33158 4278 33210
rect 4458 33158 4460 33210
rect 4214 33156 4220 33158
rect 4276 33156 4300 33158
rect 4356 33156 4380 33158
rect 4436 33156 4460 33158
rect 4516 33156 4522 33158
rect 4214 33136 4522 33156
rect 4214 32124 4522 32144
rect 4214 32122 4220 32124
rect 4276 32122 4300 32124
rect 4356 32122 4380 32124
rect 4436 32122 4460 32124
rect 4516 32122 4522 32124
rect 4276 32070 4278 32122
rect 4458 32070 4460 32122
rect 4214 32068 4220 32070
rect 4276 32068 4300 32070
rect 4356 32068 4380 32070
rect 4436 32068 4460 32070
rect 4516 32068 4522 32070
rect 4214 32048 4522 32068
rect 4214 31036 4522 31056
rect 4214 31034 4220 31036
rect 4276 31034 4300 31036
rect 4356 31034 4380 31036
rect 4436 31034 4460 31036
rect 4516 31034 4522 31036
rect 4276 30982 4278 31034
rect 4458 30982 4460 31034
rect 4214 30980 4220 30982
rect 4276 30980 4300 30982
rect 4356 30980 4380 30982
rect 4436 30980 4460 30982
rect 4516 30980 4522 30982
rect 4214 30960 4522 30980
rect 4214 29948 4522 29968
rect 4214 29946 4220 29948
rect 4276 29946 4300 29948
rect 4356 29946 4380 29948
rect 4436 29946 4460 29948
rect 4516 29946 4522 29948
rect 4276 29894 4278 29946
rect 4458 29894 4460 29946
rect 4214 29892 4220 29894
rect 4276 29892 4300 29894
rect 4356 29892 4380 29894
rect 4436 29892 4460 29894
rect 4516 29892 4522 29894
rect 4214 29872 4522 29892
rect 4214 28860 4522 28880
rect 4214 28858 4220 28860
rect 4276 28858 4300 28860
rect 4356 28858 4380 28860
rect 4436 28858 4460 28860
rect 4516 28858 4522 28860
rect 4276 28806 4278 28858
rect 4458 28806 4460 28858
rect 4214 28804 4220 28806
rect 4276 28804 4300 28806
rect 4356 28804 4380 28806
rect 4436 28804 4460 28806
rect 4516 28804 4522 28806
rect 4214 28784 4522 28804
rect 4214 27772 4522 27792
rect 4214 27770 4220 27772
rect 4276 27770 4300 27772
rect 4356 27770 4380 27772
rect 4436 27770 4460 27772
rect 4516 27770 4522 27772
rect 4276 27718 4278 27770
rect 4458 27718 4460 27770
rect 4214 27716 4220 27718
rect 4276 27716 4300 27718
rect 4356 27716 4380 27718
rect 4436 27716 4460 27718
rect 4516 27716 4522 27718
rect 4214 27696 4522 27716
rect 4214 26684 4522 26704
rect 4214 26682 4220 26684
rect 4276 26682 4300 26684
rect 4356 26682 4380 26684
rect 4436 26682 4460 26684
rect 4516 26682 4522 26684
rect 4276 26630 4278 26682
rect 4458 26630 4460 26682
rect 4214 26628 4220 26630
rect 4276 26628 4300 26630
rect 4356 26628 4380 26630
rect 4436 26628 4460 26630
rect 4516 26628 4522 26630
rect 4214 26608 4522 26628
rect 4214 25596 4522 25616
rect 4214 25594 4220 25596
rect 4276 25594 4300 25596
rect 4356 25594 4380 25596
rect 4436 25594 4460 25596
rect 4516 25594 4522 25596
rect 4276 25542 4278 25594
rect 4458 25542 4460 25594
rect 4214 25540 4220 25542
rect 4276 25540 4300 25542
rect 4356 25540 4380 25542
rect 4436 25540 4460 25542
rect 4516 25540 4522 25542
rect 4214 25520 4522 25540
rect 4214 24508 4522 24528
rect 4214 24506 4220 24508
rect 4276 24506 4300 24508
rect 4356 24506 4380 24508
rect 4436 24506 4460 24508
rect 4516 24506 4522 24508
rect 4276 24454 4278 24506
rect 4458 24454 4460 24506
rect 4214 24452 4220 24454
rect 4276 24452 4300 24454
rect 4356 24452 4380 24454
rect 4436 24452 4460 24454
rect 4516 24452 4522 24454
rect 4214 24432 4522 24452
rect 4214 23420 4522 23440
rect 4214 23418 4220 23420
rect 4276 23418 4300 23420
rect 4356 23418 4380 23420
rect 4436 23418 4460 23420
rect 4516 23418 4522 23420
rect 4276 23366 4278 23418
rect 4458 23366 4460 23418
rect 4214 23364 4220 23366
rect 4276 23364 4300 23366
rect 4356 23364 4380 23366
rect 4436 23364 4460 23366
rect 4516 23364 4522 23366
rect 4214 23344 4522 23364
rect 4214 22332 4522 22352
rect 4214 22330 4220 22332
rect 4276 22330 4300 22332
rect 4356 22330 4380 22332
rect 4436 22330 4460 22332
rect 4516 22330 4522 22332
rect 4276 22278 4278 22330
rect 4458 22278 4460 22330
rect 4214 22276 4220 22278
rect 4276 22276 4300 22278
rect 4356 22276 4380 22278
rect 4436 22276 4460 22278
rect 4516 22276 4522 22278
rect 4214 22256 4522 22276
rect 4214 21244 4522 21264
rect 4214 21242 4220 21244
rect 4276 21242 4300 21244
rect 4356 21242 4380 21244
rect 4436 21242 4460 21244
rect 4516 21242 4522 21244
rect 4276 21190 4278 21242
rect 4458 21190 4460 21242
rect 4214 21188 4220 21190
rect 4276 21188 4300 21190
rect 4356 21188 4380 21190
rect 4436 21188 4460 21190
rect 4516 21188 4522 21190
rect 4214 21168 4522 21188
rect 4214 20156 4522 20176
rect 4214 20154 4220 20156
rect 4276 20154 4300 20156
rect 4356 20154 4380 20156
rect 4436 20154 4460 20156
rect 4516 20154 4522 20156
rect 4276 20102 4278 20154
rect 4458 20102 4460 20154
rect 4214 20100 4220 20102
rect 4276 20100 4300 20102
rect 4356 20100 4380 20102
rect 4436 20100 4460 20102
rect 4516 20100 4522 20102
rect 4214 20080 4522 20100
rect 4214 19068 4522 19088
rect 4214 19066 4220 19068
rect 4276 19066 4300 19068
rect 4356 19066 4380 19068
rect 4436 19066 4460 19068
rect 4516 19066 4522 19068
rect 4276 19014 4278 19066
rect 4458 19014 4460 19066
rect 4214 19012 4220 19014
rect 4276 19012 4300 19014
rect 4356 19012 4380 19014
rect 4436 19012 4460 19014
rect 4516 19012 4522 19014
rect 4214 18992 4522 19012
rect 4214 17980 4522 18000
rect 4214 17978 4220 17980
rect 4276 17978 4300 17980
rect 4356 17978 4380 17980
rect 4436 17978 4460 17980
rect 4516 17978 4522 17980
rect 4276 17926 4278 17978
rect 4458 17926 4460 17978
rect 4214 17924 4220 17926
rect 4276 17924 4300 17926
rect 4356 17924 4380 17926
rect 4436 17924 4460 17926
rect 4516 17924 4522 17926
rect 4214 17904 4522 17924
rect 4214 16892 4522 16912
rect 4214 16890 4220 16892
rect 4276 16890 4300 16892
rect 4356 16890 4380 16892
rect 4436 16890 4460 16892
rect 4516 16890 4522 16892
rect 4276 16838 4278 16890
rect 4458 16838 4460 16890
rect 4214 16836 4220 16838
rect 4276 16836 4300 16838
rect 4356 16836 4380 16838
rect 4436 16836 4460 16838
rect 4516 16836 4522 16838
rect 4214 16816 4522 16836
rect 4632 16574 4660 35022
rect 8220 26042 8248 56238
rect 9140 55418 9168 56238
rect 25976 55826 26004 56782
rect 26056 56228 26108 56234
rect 26056 56170 26108 56176
rect 25964 55820 26016 55826
rect 25964 55762 26016 55768
rect 19574 55516 19882 55536
rect 19574 55514 19580 55516
rect 19636 55514 19660 55516
rect 19716 55514 19740 55516
rect 19796 55514 19820 55516
rect 19876 55514 19882 55516
rect 19636 55462 19638 55514
rect 19818 55462 19820 55514
rect 19574 55460 19580 55462
rect 19636 55460 19660 55462
rect 19716 55460 19740 55462
rect 19796 55460 19820 55462
rect 19876 55460 19882 55462
rect 19574 55440 19882 55460
rect 9128 55412 9180 55418
rect 9128 55354 9180 55360
rect 26068 55282 26096 56170
rect 26436 55826 26464 59200
rect 33508 56840 33560 56846
rect 33508 56782 33560 56788
rect 33520 56370 33548 56782
rect 33508 56364 33560 56370
rect 33508 56306 33560 56312
rect 34164 56302 34192 59200
rect 34934 57148 35242 57168
rect 34934 57146 34940 57148
rect 34996 57146 35020 57148
rect 35076 57146 35100 57148
rect 35156 57146 35180 57148
rect 35236 57146 35242 57148
rect 34996 57094 34998 57146
rect 35178 57094 35180 57146
rect 34934 57092 34940 57094
rect 34996 57092 35020 57094
rect 35076 57092 35100 57094
rect 35156 57092 35180 57094
rect 35236 57092 35242 57094
rect 34934 57072 35242 57092
rect 35716 56840 35768 56846
rect 35716 56782 35768 56788
rect 33692 56296 33744 56302
rect 33692 56238 33744 56244
rect 34152 56296 34204 56302
rect 34152 56238 34204 56244
rect 33704 55962 33732 56238
rect 34934 56060 35242 56080
rect 34934 56058 34940 56060
rect 34996 56058 35020 56060
rect 35076 56058 35100 56060
rect 35156 56058 35180 56060
rect 35236 56058 35242 56060
rect 34996 56006 34998 56058
rect 35178 56006 35180 56058
rect 34934 56004 34940 56006
rect 34996 56004 35020 56006
rect 35076 56004 35100 56006
rect 35156 56004 35180 56006
rect 35236 56004 35242 56006
rect 34934 55984 35242 56004
rect 33692 55956 33744 55962
rect 33692 55898 33744 55904
rect 35728 55826 35756 56782
rect 36096 55826 36124 59200
rect 41248 57458 41276 59200
rect 50294 57692 50602 57712
rect 50294 57690 50300 57692
rect 50356 57690 50380 57692
rect 50436 57690 50460 57692
rect 50516 57690 50540 57692
rect 50596 57690 50602 57692
rect 50356 57638 50358 57690
rect 50538 57638 50540 57690
rect 50294 57636 50300 57638
rect 50356 57636 50380 57638
rect 50436 57636 50460 57638
rect 50516 57636 50540 57638
rect 50596 57636 50602 57638
rect 50294 57616 50602 57636
rect 41236 57452 41288 57458
rect 41236 57394 41288 57400
rect 41696 57384 41748 57390
rect 41696 57326 41748 57332
rect 41708 55826 41736 57326
rect 42524 56840 42576 56846
rect 42524 56782 42576 56788
rect 43168 56840 43220 56846
rect 43168 56782 43220 56788
rect 49884 56840 49936 56846
rect 49884 56782 49936 56788
rect 42536 55826 42564 56782
rect 26424 55820 26476 55826
rect 26424 55762 26476 55768
rect 35716 55820 35768 55826
rect 35716 55762 35768 55768
rect 36084 55820 36136 55826
rect 36084 55762 36136 55768
rect 41696 55820 41748 55826
rect 41696 55762 41748 55768
rect 42524 55820 42576 55826
rect 42524 55762 42576 55768
rect 33600 55752 33652 55758
rect 33600 55694 33652 55700
rect 26148 55684 26200 55690
rect 26148 55626 26200 55632
rect 26160 55418 26188 55626
rect 26148 55412 26200 55418
rect 26148 55354 26200 55360
rect 9036 55276 9088 55282
rect 9036 55218 9088 55224
rect 26056 55276 26108 55282
rect 26056 55218 26108 55224
rect 8852 47048 8904 47054
rect 8852 46990 8904 46996
rect 8208 26036 8260 26042
rect 8208 25978 8260 25984
rect 8300 25900 8352 25906
rect 8300 25842 8352 25848
rect 8312 24818 8340 25842
rect 8300 24812 8352 24818
rect 8300 24754 8352 24760
rect 8312 23186 8340 24754
rect 8300 23180 8352 23186
rect 8300 23122 8352 23128
rect 7564 23112 7616 23118
rect 7564 23054 7616 23060
rect 7576 22642 7604 23054
rect 7564 22636 7616 22642
rect 7564 22578 7616 22584
rect 4632 16546 4752 16574
rect 4214 15804 4522 15824
rect 4214 15802 4220 15804
rect 4276 15802 4300 15804
rect 4356 15802 4380 15804
rect 4436 15802 4460 15804
rect 4516 15802 4522 15804
rect 4276 15750 4278 15802
rect 4458 15750 4460 15802
rect 4214 15748 4220 15750
rect 4276 15748 4300 15750
rect 4356 15748 4380 15750
rect 4436 15748 4460 15750
rect 4516 15748 4522 15750
rect 4214 15728 4522 15748
rect 4214 14716 4522 14736
rect 4214 14714 4220 14716
rect 4276 14714 4300 14716
rect 4356 14714 4380 14716
rect 4436 14714 4460 14716
rect 4516 14714 4522 14716
rect 4276 14662 4278 14714
rect 4458 14662 4460 14714
rect 4214 14660 4220 14662
rect 4276 14660 4300 14662
rect 4356 14660 4380 14662
rect 4436 14660 4460 14662
rect 4516 14660 4522 14662
rect 4214 14640 4522 14660
rect 4214 13628 4522 13648
rect 4214 13626 4220 13628
rect 4276 13626 4300 13628
rect 4356 13626 4380 13628
rect 4436 13626 4460 13628
rect 4516 13626 4522 13628
rect 4276 13574 4278 13626
rect 4458 13574 4460 13626
rect 4214 13572 4220 13574
rect 4276 13572 4300 13574
rect 4356 13572 4380 13574
rect 4436 13572 4460 13574
rect 4516 13572 4522 13574
rect 4214 13552 4522 13572
rect 4214 12540 4522 12560
rect 4214 12538 4220 12540
rect 4276 12538 4300 12540
rect 4356 12538 4380 12540
rect 4436 12538 4460 12540
rect 4516 12538 4522 12540
rect 4276 12486 4278 12538
rect 4458 12486 4460 12538
rect 4214 12484 4220 12486
rect 4276 12484 4300 12486
rect 4356 12484 4380 12486
rect 4436 12484 4460 12486
rect 4516 12484 4522 12486
rect 4214 12464 4522 12484
rect 4214 11452 4522 11472
rect 4214 11450 4220 11452
rect 4276 11450 4300 11452
rect 4356 11450 4380 11452
rect 4436 11450 4460 11452
rect 4516 11450 4522 11452
rect 4276 11398 4278 11450
rect 4458 11398 4460 11450
rect 4214 11396 4220 11398
rect 4276 11396 4300 11398
rect 4356 11396 4380 11398
rect 4436 11396 4460 11398
rect 4516 11396 4522 11398
rect 4214 11376 4522 11396
rect 2780 10600 2832 10606
rect 2780 10542 2832 10548
rect 2792 9625 2820 10542
rect 4214 10364 4522 10384
rect 4214 10362 4220 10364
rect 4276 10362 4300 10364
rect 4356 10362 4380 10364
rect 4436 10362 4460 10364
rect 4516 10362 4522 10364
rect 4276 10310 4278 10362
rect 4458 10310 4460 10362
rect 4214 10308 4220 10310
rect 4276 10308 4300 10310
rect 4356 10308 4380 10310
rect 4436 10308 4460 10310
rect 4516 10308 4522 10310
rect 4214 10288 4522 10308
rect 2778 9616 2834 9625
rect 2778 9551 2834 9560
rect 4214 9276 4522 9296
rect 4214 9274 4220 9276
rect 4276 9274 4300 9276
rect 4356 9274 4380 9276
rect 4436 9274 4460 9276
rect 4516 9274 4522 9276
rect 4276 9222 4278 9274
rect 4458 9222 4460 9274
rect 4214 9220 4220 9222
rect 4276 9220 4300 9222
rect 4356 9220 4380 9222
rect 4436 9220 4460 9222
rect 4516 9220 4522 9222
rect 4214 9200 4522 9220
rect 4214 8188 4522 8208
rect 4214 8186 4220 8188
rect 4276 8186 4300 8188
rect 4356 8186 4380 8188
rect 4436 8186 4460 8188
rect 4516 8186 4522 8188
rect 4276 8134 4278 8186
rect 4458 8134 4460 8186
rect 4214 8132 4220 8134
rect 4276 8132 4300 8134
rect 4356 8132 4380 8134
rect 4436 8132 4460 8134
rect 4516 8132 4522 8134
rect 4214 8112 4522 8132
rect 4214 7100 4522 7120
rect 4214 7098 4220 7100
rect 4276 7098 4300 7100
rect 4356 7098 4380 7100
rect 4436 7098 4460 7100
rect 4516 7098 4522 7100
rect 4276 7046 4278 7098
rect 4458 7046 4460 7098
rect 4214 7044 4220 7046
rect 4276 7044 4300 7046
rect 4356 7044 4380 7046
rect 4436 7044 4460 7046
rect 4516 7044 4522 7046
rect 4214 7024 4522 7044
rect 4214 6012 4522 6032
rect 4214 6010 4220 6012
rect 4276 6010 4300 6012
rect 4356 6010 4380 6012
rect 4436 6010 4460 6012
rect 4516 6010 4522 6012
rect 4276 5958 4278 6010
rect 4458 5958 4460 6010
rect 4214 5956 4220 5958
rect 4276 5956 4300 5958
rect 4356 5956 4380 5958
rect 4436 5956 4460 5958
rect 4516 5956 4522 5958
rect 4214 5936 4522 5956
rect 4214 4924 4522 4944
rect 4214 4922 4220 4924
rect 4276 4922 4300 4924
rect 4356 4922 4380 4924
rect 4436 4922 4460 4924
rect 4516 4922 4522 4924
rect 4276 4870 4278 4922
rect 4458 4870 4460 4922
rect 4214 4868 4220 4870
rect 4276 4868 4300 4870
rect 4356 4868 4380 4870
rect 4436 4868 4460 4870
rect 4516 4868 4522 4870
rect 2778 4856 2834 4865
rect 4214 4848 4522 4868
rect 2778 4791 2834 4800
rect 2504 4616 2556 4622
rect 2504 4558 2556 4564
rect 2136 4480 2188 4486
rect 2136 4422 2188 4428
rect 2148 4214 2176 4422
rect 2136 4208 2188 4214
rect 2136 4150 2188 4156
rect 1952 4140 2004 4146
rect 1952 4082 2004 4088
rect 2792 4078 2820 4791
rect 4724 4078 4752 16546
rect 7576 4146 7604 22578
rect 8864 22438 8892 46990
rect 9048 35086 9076 55218
rect 19574 54428 19882 54448
rect 19574 54426 19580 54428
rect 19636 54426 19660 54428
rect 19716 54426 19740 54428
rect 19796 54426 19820 54428
rect 19876 54426 19882 54428
rect 19636 54374 19638 54426
rect 19818 54374 19820 54426
rect 19574 54372 19580 54374
rect 19636 54372 19660 54374
rect 19716 54372 19740 54374
rect 19796 54372 19820 54374
rect 19876 54372 19882 54374
rect 19574 54352 19882 54372
rect 19574 53340 19882 53360
rect 19574 53338 19580 53340
rect 19636 53338 19660 53340
rect 19716 53338 19740 53340
rect 19796 53338 19820 53340
rect 19876 53338 19882 53340
rect 19636 53286 19638 53338
rect 19818 53286 19820 53338
rect 19574 53284 19580 53286
rect 19636 53284 19660 53286
rect 19716 53284 19740 53286
rect 19796 53284 19820 53286
rect 19876 53284 19882 53286
rect 19574 53264 19882 53284
rect 19574 52252 19882 52272
rect 19574 52250 19580 52252
rect 19636 52250 19660 52252
rect 19716 52250 19740 52252
rect 19796 52250 19820 52252
rect 19876 52250 19882 52252
rect 19636 52198 19638 52250
rect 19818 52198 19820 52250
rect 19574 52196 19580 52198
rect 19636 52196 19660 52198
rect 19716 52196 19740 52198
rect 19796 52196 19820 52198
rect 19876 52196 19882 52198
rect 19574 52176 19882 52196
rect 19574 51164 19882 51184
rect 19574 51162 19580 51164
rect 19636 51162 19660 51164
rect 19716 51162 19740 51164
rect 19796 51162 19820 51164
rect 19876 51162 19882 51164
rect 19636 51110 19638 51162
rect 19818 51110 19820 51162
rect 19574 51108 19580 51110
rect 19636 51108 19660 51110
rect 19716 51108 19740 51110
rect 19796 51108 19820 51110
rect 19876 51108 19882 51110
rect 19574 51088 19882 51108
rect 19574 50076 19882 50096
rect 19574 50074 19580 50076
rect 19636 50074 19660 50076
rect 19716 50074 19740 50076
rect 19796 50074 19820 50076
rect 19876 50074 19882 50076
rect 19636 50022 19638 50074
rect 19818 50022 19820 50074
rect 19574 50020 19580 50022
rect 19636 50020 19660 50022
rect 19716 50020 19740 50022
rect 19796 50020 19820 50022
rect 19876 50020 19882 50022
rect 19574 50000 19882 50020
rect 19574 48988 19882 49008
rect 19574 48986 19580 48988
rect 19636 48986 19660 48988
rect 19716 48986 19740 48988
rect 19796 48986 19820 48988
rect 19876 48986 19882 48988
rect 19636 48934 19638 48986
rect 19818 48934 19820 48986
rect 19574 48932 19580 48934
rect 19636 48932 19660 48934
rect 19716 48932 19740 48934
rect 19796 48932 19820 48934
rect 19876 48932 19882 48934
rect 19574 48912 19882 48932
rect 19574 47900 19882 47920
rect 19574 47898 19580 47900
rect 19636 47898 19660 47900
rect 19716 47898 19740 47900
rect 19796 47898 19820 47900
rect 19876 47898 19882 47900
rect 19636 47846 19638 47898
rect 19818 47846 19820 47898
rect 19574 47844 19580 47846
rect 19636 47844 19660 47846
rect 19716 47844 19740 47846
rect 19796 47844 19820 47846
rect 19876 47844 19882 47846
rect 19574 47824 19882 47844
rect 19574 46812 19882 46832
rect 19574 46810 19580 46812
rect 19636 46810 19660 46812
rect 19716 46810 19740 46812
rect 19796 46810 19820 46812
rect 19876 46810 19882 46812
rect 19636 46758 19638 46810
rect 19818 46758 19820 46810
rect 19574 46756 19580 46758
rect 19636 46756 19660 46758
rect 19716 46756 19740 46758
rect 19796 46756 19820 46758
rect 19876 46756 19882 46758
rect 19574 46736 19882 46756
rect 19574 45724 19882 45744
rect 19574 45722 19580 45724
rect 19636 45722 19660 45724
rect 19716 45722 19740 45724
rect 19796 45722 19820 45724
rect 19876 45722 19882 45724
rect 19636 45670 19638 45722
rect 19818 45670 19820 45722
rect 19574 45668 19580 45670
rect 19636 45668 19660 45670
rect 19716 45668 19740 45670
rect 19796 45668 19820 45670
rect 19876 45668 19882 45670
rect 19574 45648 19882 45668
rect 19574 44636 19882 44656
rect 19574 44634 19580 44636
rect 19636 44634 19660 44636
rect 19716 44634 19740 44636
rect 19796 44634 19820 44636
rect 19876 44634 19882 44636
rect 19636 44582 19638 44634
rect 19818 44582 19820 44634
rect 19574 44580 19580 44582
rect 19636 44580 19660 44582
rect 19716 44580 19740 44582
rect 19796 44580 19820 44582
rect 19876 44580 19882 44582
rect 19574 44560 19882 44580
rect 19574 43548 19882 43568
rect 19574 43546 19580 43548
rect 19636 43546 19660 43548
rect 19716 43546 19740 43548
rect 19796 43546 19820 43548
rect 19876 43546 19882 43548
rect 19636 43494 19638 43546
rect 19818 43494 19820 43546
rect 19574 43492 19580 43494
rect 19636 43492 19660 43494
rect 19716 43492 19740 43494
rect 19796 43492 19820 43494
rect 19876 43492 19882 43494
rect 19574 43472 19882 43492
rect 9588 42696 9640 42702
rect 9588 42638 9640 42644
rect 9600 42090 9628 42638
rect 19574 42460 19882 42480
rect 19574 42458 19580 42460
rect 19636 42458 19660 42460
rect 19716 42458 19740 42460
rect 19796 42458 19820 42460
rect 19876 42458 19882 42460
rect 19636 42406 19638 42458
rect 19818 42406 19820 42458
rect 19574 42404 19580 42406
rect 19636 42404 19660 42406
rect 19716 42404 19740 42406
rect 19796 42404 19820 42406
rect 19876 42404 19882 42406
rect 19574 42384 19882 42404
rect 33612 42090 33640 55694
rect 35900 55684 35952 55690
rect 35900 55626 35952 55632
rect 35912 55418 35940 55626
rect 35900 55412 35952 55418
rect 35900 55354 35952 55360
rect 34934 54972 35242 54992
rect 34934 54970 34940 54972
rect 34996 54970 35020 54972
rect 35076 54970 35100 54972
rect 35156 54970 35180 54972
rect 35236 54970 35242 54972
rect 34996 54918 34998 54970
rect 35178 54918 35180 54970
rect 34934 54916 34940 54918
rect 34996 54916 35020 54918
rect 35076 54916 35100 54918
rect 35156 54916 35180 54918
rect 35236 54916 35242 54918
rect 34934 54896 35242 54916
rect 41708 54738 41736 55762
rect 42708 55752 42760 55758
rect 42708 55694 42760 55700
rect 42720 55418 42748 55694
rect 42984 55616 43036 55622
rect 42984 55558 43036 55564
rect 43076 55616 43128 55622
rect 43076 55558 43128 55564
rect 42708 55412 42760 55418
rect 42708 55354 42760 55360
rect 42340 55072 42392 55078
rect 42340 55014 42392 55020
rect 42352 54738 42380 55014
rect 41696 54732 41748 54738
rect 41696 54674 41748 54680
rect 42340 54732 42392 54738
rect 42340 54674 42392 54680
rect 34934 53884 35242 53904
rect 34934 53882 34940 53884
rect 34996 53882 35020 53884
rect 35076 53882 35100 53884
rect 35156 53882 35180 53884
rect 35236 53882 35242 53884
rect 34996 53830 34998 53882
rect 35178 53830 35180 53882
rect 34934 53828 34940 53830
rect 34996 53828 35020 53830
rect 35076 53828 35100 53830
rect 35156 53828 35180 53830
rect 35236 53828 35242 53830
rect 34934 53808 35242 53828
rect 42352 53106 42380 54674
rect 42996 54534 43024 55558
rect 43088 54670 43116 55558
rect 43180 54738 43208 56782
rect 49896 56370 49924 56782
rect 50294 56604 50602 56624
rect 50294 56602 50300 56604
rect 50356 56602 50380 56604
rect 50436 56602 50460 56604
rect 50516 56602 50540 56604
rect 50596 56602 50602 56604
rect 50356 56550 50358 56602
rect 50538 56550 50540 56602
rect 50294 56548 50300 56550
rect 50356 56548 50380 56550
rect 50436 56548 50460 56550
rect 50516 56548 50540 56550
rect 50596 56548 50602 56550
rect 50294 56528 50602 56548
rect 49884 56364 49936 56370
rect 49884 56306 49936 56312
rect 50908 56302 50936 59200
rect 52840 56930 52868 59200
rect 52840 56902 52960 56930
rect 52828 56840 52880 56846
rect 52828 56782 52880 56788
rect 52840 56370 52868 56782
rect 52828 56364 52880 56370
rect 52828 56306 52880 56312
rect 44364 56296 44416 56302
rect 44364 56238 44416 56244
rect 45100 56296 45152 56302
rect 45100 56238 45152 56244
rect 50252 56296 50304 56302
rect 50252 56238 50304 56244
rect 50896 56296 50948 56302
rect 50896 56238 50948 56244
rect 43720 56160 43772 56166
rect 43720 56102 43772 56108
rect 43444 55752 43496 55758
rect 43444 55694 43496 55700
rect 43456 55282 43484 55694
rect 43536 55412 43588 55418
rect 43536 55354 43588 55360
rect 43444 55276 43496 55282
rect 43444 55218 43496 55224
rect 43168 54732 43220 54738
rect 43168 54674 43220 54680
rect 43076 54664 43128 54670
rect 43076 54606 43128 54612
rect 43548 54534 43576 55354
rect 43732 55214 43760 56102
rect 44376 55962 44404 56238
rect 44364 55956 44416 55962
rect 44364 55898 44416 55904
rect 44180 55276 44232 55282
rect 44180 55218 44232 55224
rect 43720 55208 43772 55214
rect 43720 55150 43772 55156
rect 42984 54528 43036 54534
rect 42984 54470 43036 54476
rect 43536 54528 43588 54534
rect 43536 54470 43588 54476
rect 42892 53576 42944 53582
rect 42892 53518 42944 53524
rect 42340 53100 42392 53106
rect 42340 53042 42392 53048
rect 34934 52796 35242 52816
rect 34934 52794 34940 52796
rect 34996 52794 35020 52796
rect 35076 52794 35100 52796
rect 35156 52794 35180 52796
rect 35236 52794 35242 52796
rect 34996 52742 34998 52794
rect 35178 52742 35180 52794
rect 34934 52740 34940 52742
rect 34996 52740 35020 52742
rect 35076 52740 35100 52742
rect 35156 52740 35180 52742
rect 35236 52740 35242 52742
rect 34934 52720 35242 52740
rect 42352 52578 42380 53042
rect 42904 53038 42932 53518
rect 42996 53106 43024 54470
rect 44192 53242 44220 55218
rect 45112 54874 45140 56238
rect 50264 55962 50292 56238
rect 52932 56234 52960 56902
rect 53196 56296 53248 56302
rect 53196 56238 53248 56244
rect 50344 56228 50396 56234
rect 50344 56170 50396 56176
rect 52920 56228 52972 56234
rect 52920 56170 52972 56176
rect 50252 55956 50304 55962
rect 50252 55898 50304 55904
rect 50356 55758 50384 56170
rect 53208 55962 53236 56238
rect 53196 55956 53248 55962
rect 53196 55898 53248 55904
rect 49700 55752 49752 55758
rect 49700 55694 49752 55700
rect 50344 55752 50396 55758
rect 50344 55694 50396 55700
rect 56876 55752 56928 55758
rect 56876 55694 56928 55700
rect 49712 55418 49740 55694
rect 55588 55684 55640 55690
rect 55588 55626 55640 55632
rect 50294 55516 50602 55536
rect 50294 55514 50300 55516
rect 50356 55514 50380 55516
rect 50436 55514 50460 55516
rect 50516 55514 50540 55516
rect 50596 55514 50602 55516
rect 50356 55462 50358 55514
rect 50538 55462 50540 55514
rect 50294 55460 50300 55462
rect 50356 55460 50380 55462
rect 50436 55460 50460 55462
rect 50516 55460 50540 55462
rect 50596 55460 50602 55462
rect 50294 55440 50602 55460
rect 49700 55412 49752 55418
rect 49700 55354 49752 55360
rect 45100 54868 45152 54874
rect 45100 54810 45152 54816
rect 50294 54428 50602 54448
rect 50294 54426 50300 54428
rect 50356 54426 50380 54428
rect 50436 54426 50460 54428
rect 50516 54426 50540 54428
rect 50596 54426 50602 54428
rect 50356 54374 50358 54426
rect 50538 54374 50540 54426
rect 50294 54372 50300 54374
rect 50356 54372 50380 54374
rect 50436 54372 50460 54374
rect 50516 54372 50540 54374
rect 50596 54372 50602 54374
rect 50294 54352 50602 54372
rect 46480 54188 46532 54194
rect 46480 54130 46532 54136
rect 46296 53984 46348 53990
rect 46296 53926 46348 53932
rect 45284 53712 45336 53718
rect 45284 53654 45336 53660
rect 44180 53236 44232 53242
rect 44180 53178 44232 53184
rect 42984 53100 43036 53106
rect 42984 53042 43036 53048
rect 42892 53032 42944 53038
rect 42892 52974 42944 52980
rect 42800 52692 42852 52698
rect 42800 52634 42852 52640
rect 42260 52562 42380 52578
rect 42248 52556 42380 52562
rect 42300 52550 42380 52556
rect 42248 52498 42300 52504
rect 42352 51814 42380 52550
rect 42616 52488 42668 52494
rect 42616 52430 42668 52436
rect 42628 52154 42656 52430
rect 42616 52148 42668 52154
rect 42616 52090 42668 52096
rect 42812 52018 42840 52634
rect 42996 52358 43024 53042
rect 43628 53032 43680 53038
rect 43628 52974 43680 52980
rect 43640 52698 43668 52974
rect 43628 52692 43680 52698
rect 43628 52634 43680 52640
rect 45296 52494 45324 53654
rect 45744 53576 45796 53582
rect 45744 53518 45796 53524
rect 45928 53576 45980 53582
rect 45928 53518 45980 53524
rect 45652 53440 45704 53446
rect 45652 53382 45704 53388
rect 45284 52488 45336 52494
rect 45284 52430 45336 52436
rect 42984 52352 43036 52358
rect 42984 52294 43036 52300
rect 43812 52352 43864 52358
rect 43812 52294 43864 52300
rect 43824 52154 43852 52294
rect 45664 52154 45692 53382
rect 45756 52154 45784 53518
rect 45940 52902 45968 53518
rect 46308 53174 46336 53926
rect 46492 53786 46520 54130
rect 47676 54120 47728 54126
rect 47676 54062 47728 54068
rect 46480 53780 46532 53786
rect 46480 53722 46532 53728
rect 47688 53514 47716 54062
rect 49608 53780 49660 53786
rect 49608 53722 49660 53728
rect 47676 53508 47728 53514
rect 47676 53450 47728 53456
rect 46296 53168 46348 53174
rect 46296 53110 46348 53116
rect 47688 53038 47716 53450
rect 48136 53100 48188 53106
rect 48136 53042 48188 53048
rect 48872 53100 48924 53106
rect 48872 53042 48924 53048
rect 46940 53032 46992 53038
rect 46940 52974 46992 52980
rect 47584 53032 47636 53038
rect 47584 52974 47636 52980
rect 47676 53032 47728 53038
rect 47676 52974 47728 52980
rect 45928 52896 45980 52902
rect 46952 52850 46980 52974
rect 45928 52838 45980 52844
rect 43812 52148 43864 52154
rect 43812 52090 43864 52096
rect 45652 52148 45704 52154
rect 45652 52090 45704 52096
rect 45744 52148 45796 52154
rect 45744 52090 45796 52096
rect 42800 52012 42852 52018
rect 42800 51954 42852 51960
rect 43536 51944 43588 51950
rect 43536 51886 43588 51892
rect 42340 51808 42392 51814
rect 42340 51750 42392 51756
rect 34934 51708 35242 51728
rect 34934 51706 34940 51708
rect 34996 51706 35020 51708
rect 35076 51706 35100 51708
rect 35156 51706 35180 51708
rect 35236 51706 35242 51708
rect 34996 51654 34998 51706
rect 35178 51654 35180 51706
rect 34934 51652 34940 51654
rect 34996 51652 35020 51654
rect 35076 51652 35100 51654
rect 35156 51652 35180 51654
rect 35236 51652 35242 51654
rect 34934 51632 35242 51652
rect 34934 50620 35242 50640
rect 34934 50618 34940 50620
rect 34996 50618 35020 50620
rect 35076 50618 35100 50620
rect 35156 50618 35180 50620
rect 35236 50618 35242 50620
rect 34996 50566 34998 50618
rect 35178 50566 35180 50618
rect 34934 50564 34940 50566
rect 34996 50564 35020 50566
rect 35076 50564 35100 50566
rect 35156 50564 35180 50566
rect 35236 50564 35242 50566
rect 34934 50544 35242 50564
rect 36268 50312 36320 50318
rect 36268 50254 36320 50260
rect 40500 50312 40552 50318
rect 40500 50254 40552 50260
rect 34934 49532 35242 49552
rect 34934 49530 34940 49532
rect 34996 49530 35020 49532
rect 35076 49530 35100 49532
rect 35156 49530 35180 49532
rect 35236 49530 35242 49532
rect 34996 49478 34998 49530
rect 35178 49478 35180 49530
rect 34934 49476 34940 49478
rect 34996 49476 35020 49478
rect 35076 49476 35100 49478
rect 35156 49476 35180 49478
rect 35236 49476 35242 49478
rect 34934 49456 35242 49476
rect 36280 49298 36308 50254
rect 37924 50244 37976 50250
rect 37924 50186 37976 50192
rect 37936 49978 37964 50186
rect 39488 50176 39540 50182
rect 39488 50118 39540 50124
rect 37924 49972 37976 49978
rect 37924 49914 37976 49920
rect 39500 49842 39528 50118
rect 40512 49842 40540 50254
rect 42352 49842 42380 51750
rect 38108 49836 38160 49842
rect 38108 49778 38160 49784
rect 39488 49836 39540 49842
rect 39488 49778 39540 49784
rect 40500 49836 40552 49842
rect 40500 49778 40552 49784
rect 40776 49836 40828 49842
rect 40776 49778 40828 49784
rect 42340 49836 42392 49842
rect 42340 49778 42392 49784
rect 37556 49768 37608 49774
rect 37556 49710 37608 49716
rect 36268 49292 36320 49298
rect 36268 49234 36320 49240
rect 34934 48444 35242 48464
rect 34934 48442 34940 48444
rect 34996 48442 35020 48444
rect 35076 48442 35100 48444
rect 35156 48442 35180 48444
rect 35236 48442 35242 48444
rect 34996 48390 34998 48442
rect 35178 48390 35180 48442
rect 34934 48388 34940 48390
rect 34996 48388 35020 48390
rect 35076 48388 35100 48390
rect 35156 48388 35180 48390
rect 35236 48388 35242 48390
rect 34934 48368 35242 48388
rect 34934 47356 35242 47376
rect 34934 47354 34940 47356
rect 34996 47354 35020 47356
rect 35076 47354 35100 47356
rect 35156 47354 35180 47356
rect 35236 47354 35242 47356
rect 34996 47302 34998 47354
rect 35178 47302 35180 47354
rect 34934 47300 34940 47302
rect 34996 47300 35020 47302
rect 35076 47300 35100 47302
rect 35156 47300 35180 47302
rect 35236 47300 35242 47302
rect 34934 47280 35242 47300
rect 36280 47054 36308 49234
rect 36728 49156 36780 49162
rect 36728 49098 36780 49104
rect 36740 48890 36768 49098
rect 37568 48890 37596 49710
rect 37924 49088 37976 49094
rect 37924 49030 37976 49036
rect 36728 48884 36780 48890
rect 36728 48826 36780 48832
rect 37556 48884 37608 48890
rect 37556 48826 37608 48832
rect 37936 48822 37964 49030
rect 38120 48890 38148 49778
rect 38568 49700 38620 49706
rect 38568 49642 38620 49648
rect 38108 48884 38160 48890
rect 38108 48826 38160 48832
rect 38580 48822 38608 49642
rect 39500 49434 39528 49778
rect 39856 49632 39908 49638
rect 39856 49574 39908 49580
rect 39488 49428 39540 49434
rect 39488 49370 39540 49376
rect 39868 49230 39896 49574
rect 40224 49360 40276 49366
rect 40224 49302 40276 49308
rect 39856 49224 39908 49230
rect 39856 49166 39908 49172
rect 39396 49156 39448 49162
rect 39396 49098 39448 49104
rect 39488 49156 39540 49162
rect 39488 49098 39540 49104
rect 39408 48890 39436 49098
rect 39396 48884 39448 48890
rect 39396 48826 39448 48832
rect 37924 48816 37976 48822
rect 37924 48758 37976 48764
rect 38568 48816 38620 48822
rect 38568 48758 38620 48764
rect 37832 48748 37884 48754
rect 37832 48690 37884 48696
rect 36452 48680 36504 48686
rect 36452 48622 36504 48628
rect 36464 47666 36492 48622
rect 37464 48612 37516 48618
rect 37464 48554 37516 48560
rect 37476 48346 37504 48554
rect 37556 48544 37608 48550
rect 37556 48486 37608 48492
rect 37464 48340 37516 48346
rect 37464 48282 37516 48288
rect 36728 48136 36780 48142
rect 36728 48078 36780 48084
rect 36740 47666 36768 48078
rect 37372 48000 37424 48006
rect 37372 47942 37424 47948
rect 37384 47666 37412 47942
rect 36452 47660 36504 47666
rect 36452 47602 36504 47608
rect 36728 47660 36780 47666
rect 36728 47602 36780 47608
rect 37372 47660 37424 47666
rect 37372 47602 37424 47608
rect 36360 47456 36412 47462
rect 36360 47398 36412 47404
rect 36372 47190 36400 47398
rect 36360 47184 36412 47190
rect 36360 47126 36412 47132
rect 36268 47048 36320 47054
rect 36268 46990 36320 46996
rect 34934 46268 35242 46288
rect 34934 46266 34940 46268
rect 34996 46266 35020 46268
rect 35076 46266 35100 46268
rect 35156 46266 35180 46268
rect 35236 46266 35242 46268
rect 34996 46214 34998 46266
rect 35178 46214 35180 46266
rect 34934 46212 34940 46214
rect 34996 46212 35020 46214
rect 35076 46212 35100 46214
rect 35156 46212 35180 46214
rect 35236 46212 35242 46214
rect 34934 46192 35242 46212
rect 36280 46034 36308 46990
rect 36268 46028 36320 46034
rect 36268 45970 36320 45976
rect 34934 45180 35242 45200
rect 34934 45178 34940 45180
rect 34996 45178 35020 45180
rect 35076 45178 35100 45180
rect 35156 45178 35180 45180
rect 35236 45178 35242 45180
rect 34996 45126 34998 45178
rect 35178 45126 35180 45178
rect 34934 45124 34940 45126
rect 34996 45124 35020 45126
rect 35076 45124 35100 45126
rect 35156 45124 35180 45126
rect 35236 45124 35242 45126
rect 34934 45104 35242 45124
rect 36280 44402 36308 45970
rect 36360 45960 36412 45966
rect 36464 45914 36492 47602
rect 37384 46442 37412 47602
rect 37568 47598 37596 48486
rect 37844 48142 37872 48690
rect 37832 48136 37884 48142
rect 37832 48078 37884 48084
rect 38580 48074 38608 48758
rect 39500 48754 39528 49098
rect 39672 48884 39724 48890
rect 39672 48826 39724 48832
rect 39488 48748 39540 48754
rect 39488 48690 39540 48696
rect 38844 48680 38896 48686
rect 38844 48622 38896 48628
rect 38568 48068 38620 48074
rect 38568 48010 38620 48016
rect 38580 47666 38608 48010
rect 38568 47660 38620 47666
rect 38568 47602 38620 47608
rect 37556 47592 37608 47598
rect 37556 47534 37608 47540
rect 38476 47592 38528 47598
rect 38476 47534 38528 47540
rect 38200 47456 38252 47462
rect 38200 47398 38252 47404
rect 38212 47258 38240 47398
rect 38200 47252 38252 47258
rect 38200 47194 38252 47200
rect 38488 47054 38516 47534
rect 37648 47048 37700 47054
rect 37648 46990 37700 46996
rect 38476 47048 38528 47054
rect 38476 46990 38528 46996
rect 37660 46646 37688 46990
rect 38856 46866 38884 48622
rect 39500 48550 39528 48690
rect 39488 48544 39540 48550
rect 39488 48486 39540 48492
rect 39304 48136 39356 48142
rect 39304 48078 39356 48084
rect 39316 47258 39344 48078
rect 39304 47252 39356 47258
rect 39304 47194 39356 47200
rect 39684 47054 39712 48826
rect 39868 48618 39896 49166
rect 40132 49156 40184 49162
rect 40132 49098 40184 49104
rect 39948 48680 40000 48686
rect 39948 48622 40000 48628
rect 39856 48612 39908 48618
rect 39856 48554 39908 48560
rect 39960 48142 39988 48622
rect 39948 48136 40000 48142
rect 39948 48078 40000 48084
rect 40144 47122 40172 49098
rect 40236 48822 40264 49302
rect 40316 49224 40368 49230
rect 40316 49166 40368 49172
rect 40224 48816 40276 48822
rect 40224 48758 40276 48764
rect 40236 48210 40264 48758
rect 40328 48754 40356 49166
rect 40500 49088 40552 49094
rect 40500 49030 40552 49036
rect 40512 48754 40540 49030
rect 40788 48890 40816 49778
rect 41420 49632 41472 49638
rect 41420 49574 41472 49580
rect 41432 49230 41460 49574
rect 42352 49230 42380 49778
rect 42708 49632 42760 49638
rect 42708 49574 42760 49580
rect 40868 49224 40920 49230
rect 40868 49166 40920 49172
rect 41420 49224 41472 49230
rect 41420 49166 41472 49172
rect 41604 49224 41656 49230
rect 41604 49166 41656 49172
rect 42340 49224 42392 49230
rect 42340 49166 42392 49172
rect 40776 48884 40828 48890
rect 40776 48826 40828 48832
rect 40880 48754 40908 49166
rect 41328 49088 41380 49094
rect 41328 49030 41380 49036
rect 41340 48890 41368 49030
rect 41052 48884 41104 48890
rect 41052 48826 41104 48832
rect 41328 48884 41380 48890
rect 41328 48826 41380 48832
rect 40316 48748 40368 48754
rect 40316 48690 40368 48696
rect 40500 48748 40552 48754
rect 40500 48690 40552 48696
rect 40868 48748 40920 48754
rect 40868 48690 40920 48696
rect 40224 48204 40276 48210
rect 40224 48146 40276 48152
rect 41064 47802 41092 48826
rect 41616 47802 41644 49166
rect 42352 48754 42380 49166
rect 42720 48770 42748 49574
rect 43168 49088 43220 49094
rect 43168 49030 43220 49036
rect 42340 48748 42392 48754
rect 42720 48742 42932 48770
rect 43180 48754 43208 49030
rect 42340 48690 42392 48696
rect 40316 47796 40368 47802
rect 40316 47738 40368 47744
rect 41052 47796 41104 47802
rect 41052 47738 41104 47744
rect 41604 47796 41656 47802
rect 41604 47738 41656 47744
rect 40224 47592 40276 47598
rect 40224 47534 40276 47540
rect 40132 47116 40184 47122
rect 40132 47058 40184 47064
rect 39120 47048 39172 47054
rect 39120 46990 39172 46996
rect 39672 47048 39724 47054
rect 39672 46990 39724 46996
rect 38672 46838 38884 46866
rect 37648 46640 37700 46646
rect 37648 46582 37700 46588
rect 37372 46436 37424 46442
rect 37372 46378 37424 46384
rect 36412 45908 36492 45914
rect 36360 45902 36492 45908
rect 36372 45886 36492 45902
rect 36464 44946 36492 45886
rect 37280 45892 37332 45898
rect 37280 45834 37332 45840
rect 37292 45558 37320 45834
rect 37280 45552 37332 45558
rect 37280 45494 37332 45500
rect 37384 45286 37412 46378
rect 37464 46368 37516 46374
rect 37464 46310 37516 46316
rect 37476 45490 37504 46310
rect 37660 45830 37688 46582
rect 38672 46578 38700 46838
rect 39132 46578 39160 46990
rect 38660 46572 38712 46578
rect 38660 46514 38712 46520
rect 39120 46572 39172 46578
rect 39120 46514 39172 46520
rect 38672 46034 38700 46514
rect 38660 46028 38712 46034
rect 38660 45970 38712 45976
rect 37648 45824 37700 45830
rect 37648 45766 37700 45772
rect 37660 45490 37688 45766
rect 37464 45484 37516 45490
rect 37464 45426 37516 45432
rect 37648 45484 37700 45490
rect 37648 45426 37700 45432
rect 37372 45280 37424 45286
rect 37372 45222 37424 45228
rect 36452 44940 36504 44946
rect 36452 44882 36504 44888
rect 36268 44396 36320 44402
rect 36268 44338 36320 44344
rect 34934 44092 35242 44112
rect 34934 44090 34940 44092
rect 34996 44090 35020 44092
rect 35076 44090 35100 44092
rect 35156 44090 35180 44092
rect 35236 44090 35242 44092
rect 34996 44038 34998 44090
rect 35178 44038 35180 44090
rect 34934 44036 34940 44038
rect 34996 44036 35020 44038
rect 35076 44036 35100 44038
rect 35156 44036 35180 44038
rect 35236 44036 35242 44038
rect 34934 44016 35242 44036
rect 36464 43926 36492 44882
rect 37384 44878 37412 45222
rect 39488 44940 39540 44946
rect 39488 44882 39540 44888
rect 37372 44872 37424 44878
rect 37372 44814 37424 44820
rect 37464 44872 37516 44878
rect 37464 44814 37516 44820
rect 37004 44736 37056 44742
rect 37004 44678 37056 44684
rect 37016 44470 37044 44678
rect 37004 44464 37056 44470
rect 37004 44406 37056 44412
rect 37280 44396 37332 44402
rect 37280 44338 37332 44344
rect 37292 43994 37320 44338
rect 37280 43988 37332 43994
rect 37280 43930 37332 43936
rect 36452 43920 36504 43926
rect 36452 43862 36504 43868
rect 36464 43314 36492 43862
rect 36912 43648 36964 43654
rect 36912 43590 36964 43596
rect 36452 43308 36504 43314
rect 36452 43250 36504 43256
rect 34934 43004 35242 43024
rect 34934 43002 34940 43004
rect 34996 43002 35020 43004
rect 35076 43002 35100 43004
rect 35156 43002 35180 43004
rect 35236 43002 35242 43004
rect 34996 42950 34998 43002
rect 35178 42950 35180 43002
rect 34934 42948 34940 42950
rect 34996 42948 35020 42950
rect 35076 42948 35100 42950
rect 35156 42948 35180 42950
rect 35236 42948 35242 42950
rect 34934 42928 35242 42948
rect 36924 42702 36952 43590
rect 37292 43246 37320 43930
rect 37476 43790 37504 44814
rect 38660 44736 38712 44742
rect 38660 44678 38712 44684
rect 38672 44402 38700 44678
rect 39500 44538 39528 44882
rect 39684 44538 39712 46990
rect 40236 46374 40264 47534
rect 40328 46714 40356 47738
rect 41880 47592 41932 47598
rect 41880 47534 41932 47540
rect 41892 46714 41920 47534
rect 40316 46708 40368 46714
rect 40316 46650 40368 46656
rect 41880 46708 41932 46714
rect 41880 46650 41932 46656
rect 39856 46368 39908 46374
rect 39856 46310 39908 46316
rect 40224 46368 40276 46374
rect 40224 46310 40276 46316
rect 39868 45422 39896 46310
rect 40132 46028 40184 46034
rect 40132 45970 40184 45976
rect 39856 45416 39908 45422
rect 39856 45358 39908 45364
rect 39868 44878 39896 45358
rect 39856 44872 39908 44878
rect 39856 44814 39908 44820
rect 39488 44532 39540 44538
rect 39488 44474 39540 44480
rect 39672 44532 39724 44538
rect 39672 44474 39724 44480
rect 38660 44396 38712 44402
rect 38660 44338 38712 44344
rect 37924 43920 37976 43926
rect 37924 43862 37976 43868
rect 37464 43784 37516 43790
rect 37648 43784 37700 43790
rect 37516 43744 37648 43772
rect 37464 43726 37516 43732
rect 37648 43726 37700 43732
rect 37936 43722 37964 43862
rect 38292 43784 38344 43790
rect 38292 43726 38344 43732
rect 37924 43716 37976 43722
rect 37924 43658 37976 43664
rect 37280 43240 37332 43246
rect 37280 43182 37332 43188
rect 36912 42696 36964 42702
rect 36912 42638 36964 42644
rect 37292 42634 37320 43182
rect 38304 42906 38332 43726
rect 38672 43654 38700 44338
rect 39488 44192 39540 44198
rect 39488 44134 39540 44140
rect 39500 43790 39528 44134
rect 39488 43784 39540 43790
rect 39488 43726 39540 43732
rect 38660 43648 38712 43654
rect 38660 43590 38712 43596
rect 38672 43314 38700 43590
rect 39500 43314 39528 43726
rect 38660 43308 38712 43314
rect 38660 43250 38712 43256
rect 39488 43308 39540 43314
rect 39488 43250 39540 43256
rect 38672 43110 38700 43250
rect 39868 43246 39896 44814
rect 40144 44538 40172 45970
rect 40328 45626 40356 46650
rect 42352 46510 42380 48690
rect 42904 48686 42932 48742
rect 43168 48748 43220 48754
rect 43168 48690 43220 48696
rect 42892 48680 42944 48686
rect 42892 48622 42944 48628
rect 42800 47116 42852 47122
rect 42800 47058 42852 47064
rect 41788 46504 41840 46510
rect 41788 46446 41840 46452
rect 42340 46504 42392 46510
rect 42340 46446 42392 46452
rect 41800 45626 41828 46446
rect 40316 45620 40368 45626
rect 40316 45562 40368 45568
rect 41788 45620 41840 45626
rect 41788 45562 41840 45568
rect 40328 44742 40356 45562
rect 41696 45416 41748 45422
rect 41696 45358 41748 45364
rect 41708 45082 41736 45358
rect 41696 45076 41748 45082
rect 41696 45018 41748 45024
rect 41696 44872 41748 44878
rect 41696 44814 41748 44820
rect 40316 44736 40368 44742
rect 40316 44678 40368 44684
rect 40132 44532 40184 44538
rect 40132 44474 40184 44480
rect 40328 43450 40356 44678
rect 41708 44402 41736 44814
rect 41696 44396 41748 44402
rect 41696 44338 41748 44344
rect 41512 44328 41564 44334
rect 41512 44270 41564 44276
rect 41524 43858 41552 44270
rect 41512 43852 41564 43858
rect 41512 43794 41564 43800
rect 40500 43784 40552 43790
rect 40500 43726 40552 43732
rect 40316 43444 40368 43450
rect 40316 43386 40368 43392
rect 40512 43246 40540 43726
rect 41236 43444 41288 43450
rect 41236 43386 41288 43392
rect 39856 43240 39908 43246
rect 39856 43182 39908 43188
rect 40500 43240 40552 43246
rect 40500 43182 40552 43188
rect 38660 43104 38712 43110
rect 38660 43046 38712 43052
rect 38292 42900 38344 42906
rect 38292 42842 38344 42848
rect 38672 42770 38700 43046
rect 40512 42906 40540 43182
rect 40500 42900 40552 42906
rect 40500 42842 40552 42848
rect 38660 42764 38712 42770
rect 38660 42706 38712 42712
rect 37280 42628 37332 42634
rect 37280 42570 37332 42576
rect 41248 42566 41276 43386
rect 41524 43330 41552 43794
rect 41708 43450 41736 44338
rect 42708 44328 42760 44334
rect 42812 44316 42840 47058
rect 43076 47048 43128 47054
rect 43548 47036 43576 51886
rect 43824 51074 43852 52090
rect 45664 51406 45692 52090
rect 45940 52018 45968 52838
rect 46768 52822 46980 52850
rect 46768 52698 46796 52822
rect 46756 52692 46808 52698
rect 46756 52634 46808 52640
rect 46940 52692 46992 52698
rect 46940 52634 46992 52640
rect 46848 52488 46900 52494
rect 46848 52430 46900 52436
rect 46020 52148 46072 52154
rect 46020 52090 46072 52096
rect 45928 52012 45980 52018
rect 45928 51954 45980 51960
rect 45836 51468 45888 51474
rect 45836 51410 45888 51416
rect 44732 51400 44784 51406
rect 44732 51342 44784 51348
rect 45652 51400 45704 51406
rect 45652 51342 45704 51348
rect 43732 51046 43852 51074
rect 43732 49978 43760 51046
rect 44744 50930 44772 51342
rect 45468 51264 45520 51270
rect 45468 51206 45520 51212
rect 44732 50924 44784 50930
rect 44732 50866 44784 50872
rect 43812 50720 43864 50726
rect 43812 50662 43864 50668
rect 43720 49972 43772 49978
rect 43720 49914 43772 49920
rect 43628 48884 43680 48890
rect 43732 48872 43760 49914
rect 43824 49774 43852 50662
rect 43812 49768 43864 49774
rect 43812 49710 43864 49716
rect 44180 49768 44232 49774
rect 44180 49710 44232 49716
rect 44192 48890 44220 49710
rect 45100 49632 45152 49638
rect 45100 49574 45152 49580
rect 45112 49230 45140 49574
rect 45480 49298 45508 51206
rect 45848 50930 45876 51410
rect 45940 51406 45968 51954
rect 45928 51400 45980 51406
rect 45928 51342 45980 51348
rect 46032 50930 46060 52090
rect 46664 52012 46716 52018
rect 46664 51954 46716 51960
rect 46112 51944 46164 51950
rect 46112 51886 46164 51892
rect 46124 51610 46152 51886
rect 46676 51814 46704 51954
rect 46860 51814 46888 52430
rect 46952 52018 46980 52634
rect 47596 52494 47624 52974
rect 47584 52488 47636 52494
rect 47584 52430 47636 52436
rect 46940 52012 46992 52018
rect 46940 51954 46992 51960
rect 46664 51808 46716 51814
rect 46664 51750 46716 51756
rect 46848 51808 46900 51814
rect 46848 51750 46900 51756
rect 46112 51604 46164 51610
rect 46112 51546 46164 51552
rect 46124 50998 46152 51546
rect 46860 51406 46888 51750
rect 46848 51400 46900 51406
rect 46848 51342 46900 51348
rect 46112 50992 46164 50998
rect 46112 50934 46164 50940
rect 45836 50924 45888 50930
rect 45836 50866 45888 50872
rect 46020 50924 46072 50930
rect 46020 50866 46072 50872
rect 46020 50720 46072 50726
rect 46020 50662 46072 50668
rect 45468 49292 45520 49298
rect 45468 49234 45520 49240
rect 45008 49224 45060 49230
rect 45008 49166 45060 49172
rect 45100 49224 45152 49230
rect 45100 49166 45152 49172
rect 43680 48844 43760 48872
rect 44180 48884 44232 48890
rect 43628 48826 43680 48832
rect 44180 48826 44232 48832
rect 44732 48680 44784 48686
rect 44732 48622 44784 48628
rect 44744 47734 44772 48622
rect 45020 48346 45048 49166
rect 45112 48754 45140 49166
rect 45100 48748 45152 48754
rect 45100 48690 45152 48696
rect 45008 48340 45060 48346
rect 45008 48282 45060 48288
rect 46032 48210 46060 50662
rect 47492 50176 47544 50182
rect 47492 50118 47544 50124
rect 47504 49910 47532 50118
rect 47492 49904 47544 49910
rect 47492 49846 47544 49852
rect 47596 49774 47624 52430
rect 47688 50318 47716 52974
rect 47952 52964 48004 52970
rect 47952 52906 48004 52912
rect 47768 52896 47820 52902
rect 47768 52838 47820 52844
rect 47780 52494 47808 52838
rect 47768 52488 47820 52494
rect 47768 52430 47820 52436
rect 47964 52154 47992 52906
rect 48148 52698 48176 53042
rect 48136 52692 48188 52698
rect 48136 52634 48188 52640
rect 48884 52630 48912 53042
rect 49620 52970 49648 53722
rect 50294 53340 50602 53360
rect 50294 53338 50300 53340
rect 50356 53338 50380 53340
rect 50436 53338 50460 53340
rect 50516 53338 50540 53340
rect 50596 53338 50602 53340
rect 50356 53286 50358 53338
rect 50538 53286 50540 53338
rect 50294 53284 50300 53286
rect 50356 53284 50380 53286
rect 50436 53284 50460 53286
rect 50516 53284 50540 53286
rect 50596 53284 50602 53286
rect 50294 53264 50602 53284
rect 49976 53168 50028 53174
rect 49976 53110 50028 53116
rect 49608 52964 49660 52970
rect 49608 52906 49660 52912
rect 49240 52896 49292 52902
rect 49620 52850 49648 52906
rect 49240 52838 49292 52844
rect 48872 52624 48924 52630
rect 48872 52566 48924 52572
rect 47952 52148 48004 52154
rect 47952 52090 48004 52096
rect 47964 51074 47992 52090
rect 48884 52086 48912 52566
rect 49252 52494 49280 52838
rect 49528 52822 49648 52850
rect 49240 52488 49292 52494
rect 49240 52430 49292 52436
rect 49252 52086 49280 52430
rect 49528 52426 49556 52822
rect 49608 52488 49660 52494
rect 49608 52430 49660 52436
rect 49516 52420 49568 52426
rect 49516 52362 49568 52368
rect 49528 52154 49556 52362
rect 49516 52148 49568 52154
rect 49516 52090 49568 52096
rect 48320 52080 48372 52086
rect 48320 52022 48372 52028
rect 48872 52080 48924 52086
rect 48872 52022 48924 52028
rect 49240 52080 49292 52086
rect 49240 52022 49292 52028
rect 48332 51338 48360 52022
rect 49620 52018 49648 52430
rect 49988 52426 50016 53110
rect 50344 53032 50396 53038
rect 50344 52974 50396 52980
rect 50356 52630 50384 52974
rect 50436 52896 50488 52902
rect 50436 52838 50488 52844
rect 51540 52896 51592 52902
rect 51540 52838 51592 52844
rect 50344 52624 50396 52630
rect 50344 52566 50396 52572
rect 50448 52494 50476 52838
rect 50436 52488 50488 52494
rect 50436 52430 50488 52436
rect 49976 52420 50028 52426
rect 49976 52362 50028 52368
rect 49608 52012 49660 52018
rect 49608 51954 49660 51960
rect 49988 51882 50016 52362
rect 50988 52352 51040 52358
rect 50988 52294 51040 52300
rect 50294 52252 50602 52272
rect 50294 52250 50300 52252
rect 50356 52250 50380 52252
rect 50436 52250 50460 52252
rect 50516 52250 50540 52252
rect 50596 52250 50602 52252
rect 50356 52198 50358 52250
rect 50538 52198 50540 52250
rect 50294 52196 50300 52198
rect 50356 52196 50380 52198
rect 50436 52196 50460 52198
rect 50516 52196 50540 52198
rect 50596 52196 50602 52198
rect 50294 52176 50602 52196
rect 49976 51876 50028 51882
rect 49976 51818 50028 51824
rect 49424 51808 49476 51814
rect 49424 51750 49476 51756
rect 48596 51400 48648 51406
rect 48596 51342 48648 51348
rect 48320 51332 48372 51338
rect 48320 51274 48372 51280
rect 47964 51046 48084 51074
rect 47676 50312 47728 50318
rect 47676 50254 47728 50260
rect 47584 49768 47636 49774
rect 47584 49710 47636 49716
rect 46204 49088 46256 49094
rect 46204 49030 46256 49036
rect 46848 49088 46900 49094
rect 46848 49030 46900 49036
rect 46020 48204 46072 48210
rect 46020 48146 46072 48152
rect 46216 48006 46244 49030
rect 46860 48210 46888 49030
rect 47596 48890 47624 49710
rect 47584 48884 47636 48890
rect 47584 48826 47636 48832
rect 46388 48204 46440 48210
rect 46388 48146 46440 48152
rect 46848 48204 46900 48210
rect 46848 48146 46900 48152
rect 46204 48000 46256 48006
rect 46204 47942 46256 47948
rect 44732 47728 44784 47734
rect 44732 47670 44784 47676
rect 44744 47258 44772 47670
rect 44732 47252 44784 47258
rect 44732 47194 44784 47200
rect 43628 47048 43680 47054
rect 43548 47008 43628 47036
rect 43076 46990 43128 46996
rect 43628 46990 43680 46996
rect 44364 47048 44416 47054
rect 44364 46990 44416 46996
rect 43088 46510 43116 46990
rect 44376 46714 44404 46990
rect 44456 46912 44508 46918
rect 44456 46854 44508 46860
rect 44364 46708 44416 46714
rect 44364 46650 44416 46656
rect 43076 46504 43128 46510
rect 43076 46446 43128 46452
rect 44180 46436 44232 46442
rect 44180 46378 44232 46384
rect 44192 45966 44220 46378
rect 44180 45960 44232 45966
rect 44180 45902 44232 45908
rect 43076 45824 43128 45830
rect 43076 45766 43128 45772
rect 43088 44878 43116 45766
rect 44468 45490 44496 46854
rect 44744 46034 44772 47194
rect 46216 46714 46244 47942
rect 46400 47666 46428 48146
rect 47688 47802 47716 50254
rect 48056 50250 48084 51046
rect 48608 50930 48636 51342
rect 49436 50930 49464 51750
rect 49988 51066 50016 51818
rect 50620 51808 50672 51814
rect 50620 51750 50672 51756
rect 50294 51164 50602 51184
rect 50294 51162 50300 51164
rect 50356 51162 50380 51164
rect 50436 51162 50460 51164
rect 50516 51162 50540 51164
rect 50596 51162 50602 51164
rect 50356 51110 50358 51162
rect 50538 51110 50540 51162
rect 50294 51108 50300 51110
rect 50356 51108 50380 51110
rect 50436 51108 50460 51110
rect 50516 51108 50540 51110
rect 50596 51108 50602 51110
rect 50294 51088 50602 51108
rect 49976 51060 50028 51066
rect 49976 51002 50028 51008
rect 48596 50924 48648 50930
rect 48596 50866 48648 50872
rect 49424 50924 49476 50930
rect 49424 50866 49476 50872
rect 48136 50312 48188 50318
rect 48136 50254 48188 50260
rect 48044 50244 48096 50250
rect 48044 50186 48096 50192
rect 47768 49224 47820 49230
rect 47768 49166 47820 49172
rect 47780 48686 47808 49166
rect 47768 48680 47820 48686
rect 47768 48622 47820 48628
rect 47780 48346 47808 48622
rect 48056 48618 48084 50186
rect 48148 49298 48176 50254
rect 48608 49638 48636 50866
rect 49240 50720 49292 50726
rect 49240 50662 49292 50668
rect 48596 49632 48648 49638
rect 48596 49574 48648 49580
rect 48136 49292 48188 49298
rect 48136 49234 48188 49240
rect 48044 48612 48096 48618
rect 48044 48554 48096 48560
rect 48148 48346 48176 49234
rect 48608 48822 48636 49574
rect 48964 49088 49016 49094
rect 48964 49030 49016 49036
rect 48976 48890 49004 49030
rect 48964 48884 49016 48890
rect 48964 48826 49016 48832
rect 48596 48816 48648 48822
rect 48596 48758 48648 48764
rect 49252 48686 49280 50662
rect 49988 50454 50016 51002
rect 50632 50930 50660 51750
rect 51000 51406 51028 52294
rect 51552 52018 51580 52838
rect 51540 52012 51592 52018
rect 51540 51954 51592 51960
rect 52920 51808 52972 51814
rect 52920 51750 52972 51756
rect 50988 51400 51040 51406
rect 50988 51342 51040 51348
rect 50804 51264 50856 51270
rect 50804 51206 50856 51212
rect 50620 50924 50672 50930
rect 50620 50866 50672 50872
rect 50620 50720 50672 50726
rect 50620 50662 50672 50668
rect 49976 50448 50028 50454
rect 49976 50390 50028 50396
rect 50294 50076 50602 50096
rect 50294 50074 50300 50076
rect 50356 50074 50380 50076
rect 50436 50074 50460 50076
rect 50516 50074 50540 50076
rect 50596 50074 50602 50076
rect 50356 50022 50358 50074
rect 50538 50022 50540 50074
rect 50294 50020 50300 50022
rect 50356 50020 50380 50022
rect 50436 50020 50460 50022
rect 50516 50020 50540 50022
rect 50596 50020 50602 50022
rect 50294 50000 50602 50020
rect 50160 49768 50212 49774
rect 50160 49710 50212 49716
rect 50172 49434 50200 49710
rect 50160 49428 50212 49434
rect 50160 49370 50212 49376
rect 50172 49230 50200 49370
rect 50632 49298 50660 50662
rect 50712 49972 50764 49978
rect 50712 49914 50764 49920
rect 50620 49292 50672 49298
rect 50620 49234 50672 49240
rect 50160 49224 50212 49230
rect 50160 49166 50212 49172
rect 49608 49088 49660 49094
rect 49608 49030 49660 49036
rect 50620 49088 50672 49094
rect 50724 49076 50752 49914
rect 50816 49774 50844 51206
rect 50804 49768 50856 49774
rect 50804 49710 50856 49716
rect 51080 49768 51132 49774
rect 51080 49710 51132 49716
rect 51092 49434 51120 49710
rect 50804 49428 50856 49434
rect 50804 49370 50856 49376
rect 51080 49428 51132 49434
rect 51080 49370 51132 49376
rect 50816 49094 50844 49370
rect 52932 49298 52960 51750
rect 53196 49972 53248 49978
rect 53196 49914 53248 49920
rect 53208 49298 53236 49914
rect 52644 49292 52696 49298
rect 52644 49234 52696 49240
rect 52920 49292 52972 49298
rect 52920 49234 52972 49240
rect 53196 49292 53248 49298
rect 53196 49234 53248 49240
rect 51172 49224 51224 49230
rect 51172 49166 51224 49172
rect 50672 49048 50752 49076
rect 50804 49088 50856 49094
rect 50620 49030 50672 49036
rect 50804 49030 50856 49036
rect 49240 48680 49292 48686
rect 49240 48622 49292 48628
rect 49332 48680 49384 48686
rect 49332 48622 49384 48628
rect 48412 48544 48464 48550
rect 48412 48486 48464 48492
rect 47768 48340 47820 48346
rect 47768 48282 47820 48288
rect 48136 48340 48188 48346
rect 48136 48282 48188 48288
rect 47676 47796 47728 47802
rect 47676 47738 47728 47744
rect 46388 47660 46440 47666
rect 46388 47602 46440 47608
rect 46204 46708 46256 46714
rect 46204 46650 46256 46656
rect 46216 46578 46244 46650
rect 46204 46572 46256 46578
rect 46204 46514 46256 46520
rect 47032 46504 47084 46510
rect 47032 46446 47084 46452
rect 44732 46028 44784 46034
rect 44732 45970 44784 45976
rect 45928 45892 45980 45898
rect 45928 45834 45980 45840
rect 44180 45484 44232 45490
rect 44180 45426 44232 45432
rect 44456 45484 44508 45490
rect 44456 45426 44508 45432
rect 45560 45484 45612 45490
rect 45560 45426 45612 45432
rect 43904 45280 43956 45286
rect 43904 45222 43956 45228
rect 43076 44872 43128 44878
rect 43076 44814 43128 44820
rect 42760 44288 42840 44316
rect 42708 44270 42760 44276
rect 41696 43444 41748 43450
rect 41696 43386 41748 43392
rect 41524 43302 41644 43330
rect 41512 43104 41564 43110
rect 41512 43046 41564 43052
rect 41524 42770 41552 43046
rect 41512 42764 41564 42770
rect 41512 42706 41564 42712
rect 41236 42560 41288 42566
rect 41236 42502 41288 42508
rect 9588 42084 9640 42090
rect 9588 42026 9640 42032
rect 33600 42084 33652 42090
rect 33600 42026 33652 42032
rect 9036 35080 9088 35086
rect 9036 35022 9088 35028
rect 9600 24750 9628 42026
rect 34934 41916 35242 41936
rect 34934 41914 34940 41916
rect 34996 41914 35020 41916
rect 35076 41914 35100 41916
rect 35156 41914 35180 41916
rect 35236 41914 35242 41916
rect 34996 41862 34998 41914
rect 35178 41862 35180 41914
rect 34934 41860 34940 41862
rect 34996 41860 35020 41862
rect 35076 41860 35100 41862
rect 35156 41860 35180 41862
rect 35236 41860 35242 41862
rect 34934 41840 35242 41860
rect 41616 41414 41644 43302
rect 43088 42702 43116 44814
rect 43720 44804 43772 44810
rect 43720 44746 43772 44752
rect 43732 44538 43760 44746
rect 43720 44532 43772 44538
rect 43720 44474 43772 44480
rect 43916 44402 43944 45222
rect 43904 44396 43956 44402
rect 43904 44338 43956 44344
rect 44192 44334 44220 45426
rect 44468 45286 44496 45426
rect 45468 45416 45520 45422
rect 45468 45358 45520 45364
rect 44456 45280 44508 45286
rect 44456 45222 44508 45228
rect 45480 44946 45508 45358
rect 45468 44940 45520 44946
rect 45468 44882 45520 44888
rect 44456 44736 44508 44742
rect 44456 44678 44508 44684
rect 44468 44402 44496 44678
rect 44456 44396 44508 44402
rect 44456 44338 44508 44344
rect 45376 44396 45428 44402
rect 45376 44338 45428 44344
rect 44180 44328 44232 44334
rect 44180 44270 44232 44276
rect 44192 43790 44220 44270
rect 45284 44260 45336 44266
rect 45284 44202 45336 44208
rect 45296 43790 45324 44202
rect 44180 43784 44232 43790
rect 44180 43726 44232 43732
rect 45284 43784 45336 43790
rect 45284 43726 45336 43732
rect 44192 43382 44220 43726
rect 44272 43648 44324 43654
rect 44272 43590 44324 43596
rect 44180 43376 44232 43382
rect 44180 43318 44232 43324
rect 44180 43104 44232 43110
rect 44180 43046 44232 43052
rect 43076 42696 43128 42702
rect 43076 42638 43128 42644
rect 43088 42022 43116 42638
rect 43996 42628 44048 42634
rect 43996 42570 44048 42576
rect 44008 42090 44036 42570
rect 44192 42362 44220 43046
rect 44180 42356 44232 42362
rect 44180 42298 44232 42304
rect 43996 42084 44048 42090
rect 43996 42026 44048 42032
rect 43076 42016 43128 42022
rect 43076 41958 43128 41964
rect 44192 41614 44220 42298
rect 44284 42226 44312 43590
rect 45296 43314 45324 43726
rect 45284 43308 45336 43314
rect 45284 43250 45336 43256
rect 45388 43110 45416 44338
rect 45376 43104 45428 43110
rect 45376 43046 45428 43052
rect 45388 42906 45416 43046
rect 45376 42900 45428 42906
rect 45376 42842 45428 42848
rect 45480 42362 45508 44882
rect 45572 44878 45600 45426
rect 45940 45082 45968 45834
rect 47044 45558 47072 46446
rect 47780 46374 47808 48282
rect 48424 48142 48452 48486
rect 49344 48278 49372 48622
rect 49332 48272 49384 48278
rect 49332 48214 49384 48220
rect 48412 48136 48464 48142
rect 48412 48078 48464 48084
rect 48044 46708 48096 46714
rect 48044 46650 48096 46656
rect 49424 46708 49476 46714
rect 49424 46650 49476 46656
rect 47768 46368 47820 46374
rect 47768 46310 47820 46316
rect 47780 46034 47808 46310
rect 48056 46034 48084 46650
rect 47768 46028 47820 46034
rect 47768 45970 47820 45976
rect 48044 46028 48096 46034
rect 48044 45970 48096 45976
rect 48228 46028 48280 46034
rect 48228 45970 48280 45976
rect 47124 45824 47176 45830
rect 47124 45766 47176 45772
rect 48044 45824 48096 45830
rect 48044 45766 48096 45772
rect 47032 45552 47084 45558
rect 47032 45494 47084 45500
rect 47136 45422 47164 45766
rect 47400 45484 47452 45490
rect 47400 45426 47452 45432
rect 47124 45416 47176 45422
rect 47124 45358 47176 45364
rect 46664 45280 46716 45286
rect 46664 45222 46716 45228
rect 46756 45280 46808 45286
rect 46756 45222 46808 45228
rect 46676 45082 46704 45222
rect 45928 45076 45980 45082
rect 45928 45018 45980 45024
rect 46664 45076 46716 45082
rect 46664 45018 46716 45024
rect 45560 44872 45612 44878
rect 45560 44814 45612 44820
rect 46296 44872 46348 44878
rect 46296 44814 46348 44820
rect 46572 44872 46624 44878
rect 46572 44814 46624 44820
rect 45572 43450 45600 44814
rect 46308 44402 46336 44814
rect 46296 44396 46348 44402
rect 46296 44338 46348 44344
rect 46584 43994 46612 44814
rect 46768 44266 46796 45222
rect 46940 44940 46992 44946
rect 46940 44882 46992 44888
rect 46848 44872 46900 44878
rect 46848 44814 46900 44820
rect 46860 44402 46888 44814
rect 46952 44470 46980 44882
rect 47136 44810 47164 45358
rect 47412 45082 47440 45426
rect 47400 45076 47452 45082
rect 47400 45018 47452 45024
rect 48056 44878 48084 45766
rect 47676 44872 47728 44878
rect 47676 44814 47728 44820
rect 48044 44872 48096 44878
rect 48044 44814 48096 44820
rect 47124 44804 47176 44810
rect 47124 44746 47176 44752
rect 46940 44464 46992 44470
rect 46940 44406 46992 44412
rect 46848 44396 46900 44402
rect 46848 44338 46900 44344
rect 46756 44260 46808 44266
rect 46756 44202 46808 44208
rect 46572 43988 46624 43994
rect 46572 43930 46624 43936
rect 45560 43444 45612 43450
rect 45560 43386 45612 43392
rect 45928 43444 45980 43450
rect 45928 43386 45980 43392
rect 45560 43240 45612 43246
rect 45560 43182 45612 43188
rect 45572 42770 45600 43182
rect 45560 42764 45612 42770
rect 45560 42706 45612 42712
rect 45940 42702 45968 43386
rect 46952 43246 46980 44406
rect 47688 43790 47716 44814
rect 47032 43784 47084 43790
rect 47032 43726 47084 43732
rect 47676 43784 47728 43790
rect 47676 43726 47728 43732
rect 47044 43382 47072 43726
rect 47032 43376 47084 43382
rect 47032 43318 47084 43324
rect 46940 43240 46992 43246
rect 46940 43182 46992 43188
rect 46020 42764 46072 42770
rect 46020 42706 46072 42712
rect 45836 42696 45888 42702
rect 45836 42638 45888 42644
rect 45928 42696 45980 42702
rect 45928 42638 45980 42644
rect 45560 42560 45612 42566
rect 45560 42502 45612 42508
rect 45468 42356 45520 42362
rect 45468 42298 45520 42304
rect 45572 42294 45600 42502
rect 45560 42288 45612 42294
rect 45560 42230 45612 42236
rect 44272 42220 44324 42226
rect 44272 42162 44324 42168
rect 45100 42220 45152 42226
rect 45100 42162 45152 42168
rect 45112 41818 45140 42162
rect 45100 41812 45152 41818
rect 45100 41754 45152 41760
rect 44180 41608 44232 41614
rect 44180 41550 44232 41556
rect 19574 41372 19882 41392
rect 19574 41370 19580 41372
rect 19636 41370 19660 41372
rect 19716 41370 19740 41372
rect 19796 41370 19820 41372
rect 19876 41370 19882 41372
rect 19636 41318 19638 41370
rect 19818 41318 19820 41370
rect 19574 41316 19580 41318
rect 19636 41316 19660 41318
rect 19716 41316 19740 41318
rect 19796 41316 19820 41318
rect 19876 41316 19882 41318
rect 19574 41296 19882 41316
rect 41524 41386 41644 41414
rect 34934 40828 35242 40848
rect 34934 40826 34940 40828
rect 34996 40826 35020 40828
rect 35076 40826 35100 40828
rect 35156 40826 35180 40828
rect 35236 40826 35242 40828
rect 34996 40774 34998 40826
rect 35178 40774 35180 40826
rect 34934 40772 34940 40774
rect 34996 40772 35020 40774
rect 35076 40772 35100 40774
rect 35156 40772 35180 40774
rect 35236 40772 35242 40774
rect 34934 40752 35242 40772
rect 19574 40284 19882 40304
rect 19574 40282 19580 40284
rect 19636 40282 19660 40284
rect 19716 40282 19740 40284
rect 19796 40282 19820 40284
rect 19876 40282 19882 40284
rect 19636 40230 19638 40282
rect 19818 40230 19820 40282
rect 19574 40228 19580 40230
rect 19636 40228 19660 40230
rect 19716 40228 19740 40230
rect 19796 40228 19820 40230
rect 19876 40228 19882 40230
rect 19574 40208 19882 40228
rect 34934 39740 35242 39760
rect 34934 39738 34940 39740
rect 34996 39738 35020 39740
rect 35076 39738 35100 39740
rect 35156 39738 35180 39740
rect 35236 39738 35242 39740
rect 34996 39686 34998 39738
rect 35178 39686 35180 39738
rect 34934 39684 34940 39686
rect 34996 39684 35020 39686
rect 35076 39684 35100 39686
rect 35156 39684 35180 39686
rect 35236 39684 35242 39686
rect 34934 39664 35242 39684
rect 19574 39196 19882 39216
rect 19574 39194 19580 39196
rect 19636 39194 19660 39196
rect 19716 39194 19740 39196
rect 19796 39194 19820 39196
rect 19876 39194 19882 39196
rect 19636 39142 19638 39194
rect 19818 39142 19820 39194
rect 19574 39140 19580 39142
rect 19636 39140 19660 39142
rect 19716 39140 19740 39142
rect 19796 39140 19820 39142
rect 19876 39140 19882 39142
rect 19574 39120 19882 39140
rect 34934 38652 35242 38672
rect 34934 38650 34940 38652
rect 34996 38650 35020 38652
rect 35076 38650 35100 38652
rect 35156 38650 35180 38652
rect 35236 38650 35242 38652
rect 34996 38598 34998 38650
rect 35178 38598 35180 38650
rect 34934 38596 34940 38598
rect 34996 38596 35020 38598
rect 35076 38596 35100 38598
rect 35156 38596 35180 38598
rect 35236 38596 35242 38598
rect 34934 38576 35242 38596
rect 19574 38108 19882 38128
rect 19574 38106 19580 38108
rect 19636 38106 19660 38108
rect 19716 38106 19740 38108
rect 19796 38106 19820 38108
rect 19876 38106 19882 38108
rect 19636 38054 19638 38106
rect 19818 38054 19820 38106
rect 19574 38052 19580 38054
rect 19636 38052 19660 38054
rect 19716 38052 19740 38054
rect 19796 38052 19820 38054
rect 19876 38052 19882 38054
rect 19574 38032 19882 38052
rect 34934 37564 35242 37584
rect 34934 37562 34940 37564
rect 34996 37562 35020 37564
rect 35076 37562 35100 37564
rect 35156 37562 35180 37564
rect 35236 37562 35242 37564
rect 34996 37510 34998 37562
rect 35178 37510 35180 37562
rect 34934 37508 34940 37510
rect 34996 37508 35020 37510
rect 35076 37508 35100 37510
rect 35156 37508 35180 37510
rect 35236 37508 35242 37510
rect 34934 37488 35242 37508
rect 19574 37020 19882 37040
rect 19574 37018 19580 37020
rect 19636 37018 19660 37020
rect 19716 37018 19740 37020
rect 19796 37018 19820 37020
rect 19876 37018 19882 37020
rect 19636 36966 19638 37018
rect 19818 36966 19820 37018
rect 19574 36964 19580 36966
rect 19636 36964 19660 36966
rect 19716 36964 19740 36966
rect 19796 36964 19820 36966
rect 19876 36964 19882 36966
rect 19574 36944 19882 36964
rect 34934 36476 35242 36496
rect 34934 36474 34940 36476
rect 34996 36474 35020 36476
rect 35076 36474 35100 36476
rect 35156 36474 35180 36476
rect 35236 36474 35242 36476
rect 34996 36422 34998 36474
rect 35178 36422 35180 36474
rect 34934 36420 34940 36422
rect 34996 36420 35020 36422
rect 35076 36420 35100 36422
rect 35156 36420 35180 36422
rect 35236 36420 35242 36422
rect 34934 36400 35242 36420
rect 19574 35932 19882 35952
rect 19574 35930 19580 35932
rect 19636 35930 19660 35932
rect 19716 35930 19740 35932
rect 19796 35930 19820 35932
rect 19876 35930 19882 35932
rect 19636 35878 19638 35930
rect 19818 35878 19820 35930
rect 19574 35876 19580 35878
rect 19636 35876 19660 35878
rect 19716 35876 19740 35878
rect 19796 35876 19820 35878
rect 19876 35876 19882 35878
rect 19574 35856 19882 35876
rect 34934 35388 35242 35408
rect 34934 35386 34940 35388
rect 34996 35386 35020 35388
rect 35076 35386 35100 35388
rect 35156 35386 35180 35388
rect 35236 35386 35242 35388
rect 34996 35334 34998 35386
rect 35178 35334 35180 35386
rect 34934 35332 34940 35334
rect 34996 35332 35020 35334
rect 35076 35332 35100 35334
rect 35156 35332 35180 35334
rect 35236 35332 35242 35334
rect 34934 35312 35242 35332
rect 19574 34844 19882 34864
rect 19574 34842 19580 34844
rect 19636 34842 19660 34844
rect 19716 34842 19740 34844
rect 19796 34842 19820 34844
rect 19876 34842 19882 34844
rect 19636 34790 19638 34842
rect 19818 34790 19820 34842
rect 19574 34788 19580 34790
rect 19636 34788 19660 34790
rect 19716 34788 19740 34790
rect 19796 34788 19820 34790
rect 19876 34788 19882 34790
rect 19574 34768 19882 34788
rect 34934 34300 35242 34320
rect 34934 34298 34940 34300
rect 34996 34298 35020 34300
rect 35076 34298 35100 34300
rect 35156 34298 35180 34300
rect 35236 34298 35242 34300
rect 34996 34246 34998 34298
rect 35178 34246 35180 34298
rect 34934 34244 34940 34246
rect 34996 34244 35020 34246
rect 35076 34244 35100 34246
rect 35156 34244 35180 34246
rect 35236 34244 35242 34246
rect 34934 34224 35242 34244
rect 19574 33756 19882 33776
rect 19574 33754 19580 33756
rect 19636 33754 19660 33756
rect 19716 33754 19740 33756
rect 19796 33754 19820 33756
rect 19876 33754 19882 33756
rect 19636 33702 19638 33754
rect 19818 33702 19820 33754
rect 19574 33700 19580 33702
rect 19636 33700 19660 33702
rect 19716 33700 19740 33702
rect 19796 33700 19820 33702
rect 19876 33700 19882 33702
rect 19574 33680 19882 33700
rect 34934 33212 35242 33232
rect 34934 33210 34940 33212
rect 34996 33210 35020 33212
rect 35076 33210 35100 33212
rect 35156 33210 35180 33212
rect 35236 33210 35242 33212
rect 34996 33158 34998 33210
rect 35178 33158 35180 33210
rect 34934 33156 34940 33158
rect 34996 33156 35020 33158
rect 35076 33156 35100 33158
rect 35156 33156 35180 33158
rect 35236 33156 35242 33158
rect 34934 33136 35242 33156
rect 19574 32668 19882 32688
rect 19574 32666 19580 32668
rect 19636 32666 19660 32668
rect 19716 32666 19740 32668
rect 19796 32666 19820 32668
rect 19876 32666 19882 32668
rect 19636 32614 19638 32666
rect 19818 32614 19820 32666
rect 19574 32612 19580 32614
rect 19636 32612 19660 32614
rect 19716 32612 19740 32614
rect 19796 32612 19820 32614
rect 19876 32612 19882 32614
rect 19574 32592 19882 32612
rect 34934 32124 35242 32144
rect 34934 32122 34940 32124
rect 34996 32122 35020 32124
rect 35076 32122 35100 32124
rect 35156 32122 35180 32124
rect 35236 32122 35242 32124
rect 34996 32070 34998 32122
rect 35178 32070 35180 32122
rect 34934 32068 34940 32070
rect 34996 32068 35020 32070
rect 35076 32068 35100 32070
rect 35156 32068 35180 32070
rect 35236 32068 35242 32070
rect 34934 32048 35242 32068
rect 19574 31580 19882 31600
rect 19574 31578 19580 31580
rect 19636 31578 19660 31580
rect 19716 31578 19740 31580
rect 19796 31578 19820 31580
rect 19876 31578 19882 31580
rect 19636 31526 19638 31578
rect 19818 31526 19820 31578
rect 19574 31524 19580 31526
rect 19636 31524 19660 31526
rect 19716 31524 19740 31526
rect 19796 31524 19820 31526
rect 19876 31524 19882 31526
rect 19574 31504 19882 31524
rect 34934 31036 35242 31056
rect 34934 31034 34940 31036
rect 34996 31034 35020 31036
rect 35076 31034 35100 31036
rect 35156 31034 35180 31036
rect 35236 31034 35242 31036
rect 34996 30982 34998 31034
rect 35178 30982 35180 31034
rect 34934 30980 34940 30982
rect 34996 30980 35020 30982
rect 35076 30980 35100 30982
rect 35156 30980 35180 30982
rect 35236 30980 35242 30982
rect 34934 30960 35242 30980
rect 19574 30492 19882 30512
rect 19574 30490 19580 30492
rect 19636 30490 19660 30492
rect 19716 30490 19740 30492
rect 19796 30490 19820 30492
rect 19876 30490 19882 30492
rect 19636 30438 19638 30490
rect 19818 30438 19820 30490
rect 19574 30436 19580 30438
rect 19636 30436 19660 30438
rect 19716 30436 19740 30438
rect 19796 30436 19820 30438
rect 19876 30436 19882 30438
rect 19574 30416 19882 30436
rect 34934 29948 35242 29968
rect 34934 29946 34940 29948
rect 34996 29946 35020 29948
rect 35076 29946 35100 29948
rect 35156 29946 35180 29948
rect 35236 29946 35242 29948
rect 34996 29894 34998 29946
rect 35178 29894 35180 29946
rect 34934 29892 34940 29894
rect 34996 29892 35020 29894
rect 35076 29892 35100 29894
rect 35156 29892 35180 29894
rect 35236 29892 35242 29894
rect 34934 29872 35242 29892
rect 19574 29404 19882 29424
rect 19574 29402 19580 29404
rect 19636 29402 19660 29404
rect 19716 29402 19740 29404
rect 19796 29402 19820 29404
rect 19876 29402 19882 29404
rect 19636 29350 19638 29402
rect 19818 29350 19820 29402
rect 19574 29348 19580 29350
rect 19636 29348 19660 29350
rect 19716 29348 19740 29350
rect 19796 29348 19820 29350
rect 19876 29348 19882 29350
rect 19574 29328 19882 29348
rect 34934 28860 35242 28880
rect 34934 28858 34940 28860
rect 34996 28858 35020 28860
rect 35076 28858 35100 28860
rect 35156 28858 35180 28860
rect 35236 28858 35242 28860
rect 34996 28806 34998 28858
rect 35178 28806 35180 28858
rect 34934 28804 34940 28806
rect 34996 28804 35020 28806
rect 35076 28804 35100 28806
rect 35156 28804 35180 28806
rect 35236 28804 35242 28806
rect 34934 28784 35242 28804
rect 19574 28316 19882 28336
rect 19574 28314 19580 28316
rect 19636 28314 19660 28316
rect 19716 28314 19740 28316
rect 19796 28314 19820 28316
rect 19876 28314 19882 28316
rect 19636 28262 19638 28314
rect 19818 28262 19820 28314
rect 19574 28260 19580 28262
rect 19636 28260 19660 28262
rect 19716 28260 19740 28262
rect 19796 28260 19820 28262
rect 19876 28260 19882 28262
rect 19574 28240 19882 28260
rect 34934 27772 35242 27792
rect 34934 27770 34940 27772
rect 34996 27770 35020 27772
rect 35076 27770 35100 27772
rect 35156 27770 35180 27772
rect 35236 27770 35242 27772
rect 34996 27718 34998 27770
rect 35178 27718 35180 27770
rect 34934 27716 34940 27718
rect 34996 27716 35020 27718
rect 35076 27716 35100 27718
rect 35156 27716 35180 27718
rect 35236 27716 35242 27718
rect 34934 27696 35242 27716
rect 19574 27228 19882 27248
rect 19574 27226 19580 27228
rect 19636 27226 19660 27228
rect 19716 27226 19740 27228
rect 19796 27226 19820 27228
rect 19876 27226 19882 27228
rect 19636 27174 19638 27226
rect 19818 27174 19820 27226
rect 19574 27172 19580 27174
rect 19636 27172 19660 27174
rect 19716 27172 19740 27174
rect 19796 27172 19820 27174
rect 19876 27172 19882 27174
rect 19574 27152 19882 27172
rect 34934 26684 35242 26704
rect 34934 26682 34940 26684
rect 34996 26682 35020 26684
rect 35076 26682 35100 26684
rect 35156 26682 35180 26684
rect 35236 26682 35242 26684
rect 34996 26630 34998 26682
rect 35178 26630 35180 26682
rect 34934 26628 34940 26630
rect 34996 26628 35020 26630
rect 35076 26628 35100 26630
rect 35156 26628 35180 26630
rect 35236 26628 35242 26630
rect 34934 26608 35242 26628
rect 19574 26140 19882 26160
rect 19574 26138 19580 26140
rect 19636 26138 19660 26140
rect 19716 26138 19740 26140
rect 19796 26138 19820 26140
rect 19876 26138 19882 26140
rect 19636 26086 19638 26138
rect 19818 26086 19820 26138
rect 19574 26084 19580 26086
rect 19636 26084 19660 26086
rect 19716 26084 19740 26086
rect 19796 26084 19820 26086
rect 19876 26084 19882 26086
rect 19574 26064 19882 26084
rect 34934 25596 35242 25616
rect 34934 25594 34940 25596
rect 34996 25594 35020 25596
rect 35076 25594 35100 25596
rect 35156 25594 35180 25596
rect 35236 25594 35242 25596
rect 34996 25542 34998 25594
rect 35178 25542 35180 25594
rect 34934 25540 34940 25542
rect 34996 25540 35020 25542
rect 35076 25540 35100 25542
rect 35156 25540 35180 25542
rect 35236 25540 35242 25542
rect 34934 25520 35242 25540
rect 19574 25052 19882 25072
rect 19574 25050 19580 25052
rect 19636 25050 19660 25052
rect 19716 25050 19740 25052
rect 19796 25050 19820 25052
rect 19876 25050 19882 25052
rect 19636 24998 19638 25050
rect 19818 24998 19820 25050
rect 19574 24996 19580 24998
rect 19636 24996 19660 24998
rect 19716 24996 19740 24998
rect 19796 24996 19820 24998
rect 19876 24996 19882 24998
rect 19574 24976 19882 24996
rect 9588 24744 9640 24750
rect 9588 24686 9640 24692
rect 34934 24508 35242 24528
rect 34934 24506 34940 24508
rect 34996 24506 35020 24508
rect 35076 24506 35100 24508
rect 35156 24506 35180 24508
rect 35236 24506 35242 24508
rect 34996 24454 34998 24506
rect 35178 24454 35180 24506
rect 34934 24452 34940 24454
rect 34996 24452 35020 24454
rect 35076 24452 35100 24454
rect 35156 24452 35180 24454
rect 35236 24452 35242 24454
rect 34934 24432 35242 24452
rect 19574 23964 19882 23984
rect 19574 23962 19580 23964
rect 19636 23962 19660 23964
rect 19716 23962 19740 23964
rect 19796 23962 19820 23964
rect 19876 23962 19882 23964
rect 19636 23910 19638 23962
rect 19818 23910 19820 23962
rect 19574 23908 19580 23910
rect 19636 23908 19660 23910
rect 19716 23908 19740 23910
rect 19796 23908 19820 23910
rect 19876 23908 19882 23910
rect 19574 23888 19882 23908
rect 34934 23420 35242 23440
rect 34934 23418 34940 23420
rect 34996 23418 35020 23420
rect 35076 23418 35100 23420
rect 35156 23418 35180 23420
rect 35236 23418 35242 23420
rect 34996 23366 34998 23418
rect 35178 23366 35180 23418
rect 34934 23364 34940 23366
rect 34996 23364 35020 23366
rect 35076 23364 35100 23366
rect 35156 23364 35180 23366
rect 35236 23364 35242 23366
rect 34934 23344 35242 23364
rect 19574 22876 19882 22896
rect 19574 22874 19580 22876
rect 19636 22874 19660 22876
rect 19716 22874 19740 22876
rect 19796 22874 19820 22876
rect 19876 22874 19882 22876
rect 19636 22822 19638 22874
rect 19818 22822 19820 22874
rect 19574 22820 19580 22822
rect 19636 22820 19660 22822
rect 19716 22820 19740 22822
rect 19796 22820 19820 22822
rect 19876 22820 19882 22822
rect 19574 22800 19882 22820
rect 8852 22432 8904 22438
rect 8852 22374 8904 22380
rect 8864 11150 8892 22374
rect 34934 22332 35242 22352
rect 34934 22330 34940 22332
rect 34996 22330 35020 22332
rect 35076 22330 35100 22332
rect 35156 22330 35180 22332
rect 35236 22330 35242 22332
rect 34996 22278 34998 22330
rect 35178 22278 35180 22330
rect 34934 22276 34940 22278
rect 34996 22276 35020 22278
rect 35076 22276 35100 22278
rect 35156 22276 35180 22278
rect 35236 22276 35242 22278
rect 34934 22256 35242 22276
rect 19574 21788 19882 21808
rect 19574 21786 19580 21788
rect 19636 21786 19660 21788
rect 19716 21786 19740 21788
rect 19796 21786 19820 21788
rect 19876 21786 19882 21788
rect 19636 21734 19638 21786
rect 19818 21734 19820 21786
rect 19574 21732 19580 21734
rect 19636 21732 19660 21734
rect 19716 21732 19740 21734
rect 19796 21732 19820 21734
rect 19876 21732 19882 21734
rect 19574 21712 19882 21732
rect 34934 21244 35242 21264
rect 34934 21242 34940 21244
rect 34996 21242 35020 21244
rect 35076 21242 35100 21244
rect 35156 21242 35180 21244
rect 35236 21242 35242 21244
rect 34996 21190 34998 21242
rect 35178 21190 35180 21242
rect 34934 21188 34940 21190
rect 34996 21188 35020 21190
rect 35076 21188 35100 21190
rect 35156 21188 35180 21190
rect 35236 21188 35242 21190
rect 34934 21168 35242 21188
rect 19574 20700 19882 20720
rect 19574 20698 19580 20700
rect 19636 20698 19660 20700
rect 19716 20698 19740 20700
rect 19796 20698 19820 20700
rect 19876 20698 19882 20700
rect 19636 20646 19638 20698
rect 19818 20646 19820 20698
rect 19574 20644 19580 20646
rect 19636 20644 19660 20646
rect 19716 20644 19740 20646
rect 19796 20644 19820 20646
rect 19876 20644 19882 20646
rect 19574 20624 19882 20644
rect 34934 20156 35242 20176
rect 34934 20154 34940 20156
rect 34996 20154 35020 20156
rect 35076 20154 35100 20156
rect 35156 20154 35180 20156
rect 35236 20154 35242 20156
rect 34996 20102 34998 20154
rect 35178 20102 35180 20154
rect 34934 20100 34940 20102
rect 34996 20100 35020 20102
rect 35076 20100 35100 20102
rect 35156 20100 35180 20102
rect 35236 20100 35242 20102
rect 34934 20080 35242 20100
rect 19574 19612 19882 19632
rect 19574 19610 19580 19612
rect 19636 19610 19660 19612
rect 19716 19610 19740 19612
rect 19796 19610 19820 19612
rect 19876 19610 19882 19612
rect 19636 19558 19638 19610
rect 19818 19558 19820 19610
rect 19574 19556 19580 19558
rect 19636 19556 19660 19558
rect 19716 19556 19740 19558
rect 19796 19556 19820 19558
rect 19876 19556 19882 19558
rect 19574 19536 19882 19556
rect 34934 19068 35242 19088
rect 34934 19066 34940 19068
rect 34996 19066 35020 19068
rect 35076 19066 35100 19068
rect 35156 19066 35180 19068
rect 35236 19066 35242 19068
rect 34996 19014 34998 19066
rect 35178 19014 35180 19066
rect 34934 19012 34940 19014
rect 34996 19012 35020 19014
rect 35076 19012 35100 19014
rect 35156 19012 35180 19014
rect 35236 19012 35242 19014
rect 34934 18992 35242 19012
rect 19574 18524 19882 18544
rect 19574 18522 19580 18524
rect 19636 18522 19660 18524
rect 19716 18522 19740 18524
rect 19796 18522 19820 18524
rect 19876 18522 19882 18524
rect 19636 18470 19638 18522
rect 19818 18470 19820 18522
rect 19574 18468 19580 18470
rect 19636 18468 19660 18470
rect 19716 18468 19740 18470
rect 19796 18468 19820 18470
rect 19876 18468 19882 18470
rect 19574 18448 19882 18468
rect 34934 17980 35242 18000
rect 34934 17978 34940 17980
rect 34996 17978 35020 17980
rect 35076 17978 35100 17980
rect 35156 17978 35180 17980
rect 35236 17978 35242 17980
rect 34996 17926 34998 17978
rect 35178 17926 35180 17978
rect 34934 17924 34940 17926
rect 34996 17924 35020 17926
rect 35076 17924 35100 17926
rect 35156 17924 35180 17926
rect 35236 17924 35242 17926
rect 34934 17904 35242 17924
rect 19574 17436 19882 17456
rect 19574 17434 19580 17436
rect 19636 17434 19660 17436
rect 19716 17434 19740 17436
rect 19796 17434 19820 17436
rect 19876 17434 19882 17436
rect 19636 17382 19638 17434
rect 19818 17382 19820 17434
rect 19574 17380 19580 17382
rect 19636 17380 19660 17382
rect 19716 17380 19740 17382
rect 19796 17380 19820 17382
rect 19876 17380 19882 17382
rect 19574 17360 19882 17380
rect 34934 16892 35242 16912
rect 34934 16890 34940 16892
rect 34996 16890 35020 16892
rect 35076 16890 35100 16892
rect 35156 16890 35180 16892
rect 35236 16890 35242 16892
rect 34996 16838 34998 16890
rect 35178 16838 35180 16890
rect 34934 16836 34940 16838
rect 34996 16836 35020 16838
rect 35076 16836 35100 16838
rect 35156 16836 35180 16838
rect 35236 16836 35242 16838
rect 34934 16816 35242 16836
rect 19574 16348 19882 16368
rect 19574 16346 19580 16348
rect 19636 16346 19660 16348
rect 19716 16346 19740 16348
rect 19796 16346 19820 16348
rect 19876 16346 19882 16348
rect 19636 16294 19638 16346
rect 19818 16294 19820 16346
rect 19574 16292 19580 16294
rect 19636 16292 19660 16294
rect 19716 16292 19740 16294
rect 19796 16292 19820 16294
rect 19876 16292 19882 16294
rect 19574 16272 19882 16292
rect 34934 15804 35242 15824
rect 34934 15802 34940 15804
rect 34996 15802 35020 15804
rect 35076 15802 35100 15804
rect 35156 15802 35180 15804
rect 35236 15802 35242 15804
rect 34996 15750 34998 15802
rect 35178 15750 35180 15802
rect 34934 15748 34940 15750
rect 34996 15748 35020 15750
rect 35076 15748 35100 15750
rect 35156 15748 35180 15750
rect 35236 15748 35242 15750
rect 34934 15728 35242 15748
rect 19574 15260 19882 15280
rect 19574 15258 19580 15260
rect 19636 15258 19660 15260
rect 19716 15258 19740 15260
rect 19796 15258 19820 15260
rect 19876 15258 19882 15260
rect 19636 15206 19638 15258
rect 19818 15206 19820 15258
rect 19574 15204 19580 15206
rect 19636 15204 19660 15206
rect 19716 15204 19740 15206
rect 19796 15204 19820 15206
rect 19876 15204 19882 15206
rect 19574 15184 19882 15204
rect 34934 14716 35242 14736
rect 34934 14714 34940 14716
rect 34996 14714 35020 14716
rect 35076 14714 35100 14716
rect 35156 14714 35180 14716
rect 35236 14714 35242 14716
rect 34996 14662 34998 14714
rect 35178 14662 35180 14714
rect 34934 14660 34940 14662
rect 34996 14660 35020 14662
rect 35076 14660 35100 14662
rect 35156 14660 35180 14662
rect 35236 14660 35242 14662
rect 34934 14640 35242 14660
rect 19574 14172 19882 14192
rect 19574 14170 19580 14172
rect 19636 14170 19660 14172
rect 19716 14170 19740 14172
rect 19796 14170 19820 14172
rect 19876 14170 19882 14172
rect 19636 14118 19638 14170
rect 19818 14118 19820 14170
rect 19574 14116 19580 14118
rect 19636 14116 19660 14118
rect 19716 14116 19740 14118
rect 19796 14116 19820 14118
rect 19876 14116 19882 14118
rect 19574 14096 19882 14116
rect 34934 13628 35242 13648
rect 34934 13626 34940 13628
rect 34996 13626 35020 13628
rect 35076 13626 35100 13628
rect 35156 13626 35180 13628
rect 35236 13626 35242 13628
rect 34996 13574 34998 13626
rect 35178 13574 35180 13626
rect 34934 13572 34940 13574
rect 34996 13572 35020 13574
rect 35076 13572 35100 13574
rect 35156 13572 35180 13574
rect 35236 13572 35242 13574
rect 34934 13552 35242 13572
rect 19574 13084 19882 13104
rect 19574 13082 19580 13084
rect 19636 13082 19660 13084
rect 19716 13082 19740 13084
rect 19796 13082 19820 13084
rect 19876 13082 19882 13084
rect 19636 13030 19638 13082
rect 19818 13030 19820 13082
rect 19574 13028 19580 13030
rect 19636 13028 19660 13030
rect 19716 13028 19740 13030
rect 19796 13028 19820 13030
rect 19876 13028 19882 13030
rect 19574 13008 19882 13028
rect 34934 12540 35242 12560
rect 34934 12538 34940 12540
rect 34996 12538 35020 12540
rect 35076 12538 35100 12540
rect 35156 12538 35180 12540
rect 35236 12538 35242 12540
rect 34996 12486 34998 12538
rect 35178 12486 35180 12538
rect 34934 12484 34940 12486
rect 34996 12484 35020 12486
rect 35076 12484 35100 12486
rect 35156 12484 35180 12486
rect 35236 12484 35242 12486
rect 34934 12464 35242 12484
rect 19574 11996 19882 12016
rect 19574 11994 19580 11996
rect 19636 11994 19660 11996
rect 19716 11994 19740 11996
rect 19796 11994 19820 11996
rect 19876 11994 19882 11996
rect 19636 11942 19638 11994
rect 19818 11942 19820 11994
rect 19574 11940 19580 11942
rect 19636 11940 19660 11942
rect 19716 11940 19740 11942
rect 19796 11940 19820 11942
rect 19876 11940 19882 11942
rect 19574 11920 19882 11940
rect 34934 11452 35242 11472
rect 34934 11450 34940 11452
rect 34996 11450 35020 11452
rect 35076 11450 35100 11452
rect 35156 11450 35180 11452
rect 35236 11450 35242 11452
rect 34996 11398 34998 11450
rect 35178 11398 35180 11450
rect 34934 11396 34940 11398
rect 34996 11396 35020 11398
rect 35076 11396 35100 11398
rect 35156 11396 35180 11398
rect 35236 11396 35242 11398
rect 34934 11376 35242 11396
rect 8852 11144 8904 11150
rect 8852 11086 8904 11092
rect 19574 10908 19882 10928
rect 19574 10906 19580 10908
rect 19636 10906 19660 10908
rect 19716 10906 19740 10908
rect 19796 10906 19820 10908
rect 19876 10906 19882 10908
rect 19636 10854 19638 10906
rect 19818 10854 19820 10906
rect 19574 10852 19580 10854
rect 19636 10852 19660 10854
rect 19716 10852 19740 10854
rect 19796 10852 19820 10854
rect 19876 10852 19882 10854
rect 19574 10832 19882 10852
rect 34934 10364 35242 10384
rect 34934 10362 34940 10364
rect 34996 10362 35020 10364
rect 35076 10362 35100 10364
rect 35156 10362 35180 10364
rect 35236 10362 35242 10364
rect 34996 10310 34998 10362
rect 35178 10310 35180 10362
rect 34934 10308 34940 10310
rect 34996 10308 35020 10310
rect 35076 10308 35100 10310
rect 35156 10308 35180 10310
rect 35236 10308 35242 10310
rect 34934 10288 35242 10308
rect 19574 9820 19882 9840
rect 19574 9818 19580 9820
rect 19636 9818 19660 9820
rect 19716 9818 19740 9820
rect 19796 9818 19820 9820
rect 19876 9818 19882 9820
rect 19636 9766 19638 9818
rect 19818 9766 19820 9818
rect 19574 9764 19580 9766
rect 19636 9764 19660 9766
rect 19716 9764 19740 9766
rect 19796 9764 19820 9766
rect 19876 9764 19882 9766
rect 19574 9744 19882 9764
rect 34934 9276 35242 9296
rect 34934 9274 34940 9276
rect 34996 9274 35020 9276
rect 35076 9274 35100 9276
rect 35156 9274 35180 9276
rect 35236 9274 35242 9276
rect 34996 9222 34998 9274
rect 35178 9222 35180 9274
rect 34934 9220 34940 9222
rect 34996 9220 35020 9222
rect 35076 9220 35100 9222
rect 35156 9220 35180 9222
rect 35236 9220 35242 9222
rect 34934 9200 35242 9220
rect 19574 8732 19882 8752
rect 19574 8730 19580 8732
rect 19636 8730 19660 8732
rect 19716 8730 19740 8732
rect 19796 8730 19820 8732
rect 19876 8730 19882 8732
rect 19636 8678 19638 8730
rect 19818 8678 19820 8730
rect 19574 8676 19580 8678
rect 19636 8676 19660 8678
rect 19716 8676 19740 8678
rect 19796 8676 19820 8678
rect 19876 8676 19882 8678
rect 19574 8656 19882 8676
rect 34934 8188 35242 8208
rect 34934 8186 34940 8188
rect 34996 8186 35020 8188
rect 35076 8186 35100 8188
rect 35156 8186 35180 8188
rect 35236 8186 35242 8188
rect 34996 8134 34998 8186
rect 35178 8134 35180 8186
rect 34934 8132 34940 8134
rect 34996 8132 35020 8134
rect 35076 8132 35100 8134
rect 35156 8132 35180 8134
rect 35236 8132 35242 8134
rect 34934 8112 35242 8132
rect 19574 7644 19882 7664
rect 19574 7642 19580 7644
rect 19636 7642 19660 7644
rect 19716 7642 19740 7644
rect 19796 7642 19820 7644
rect 19876 7642 19882 7644
rect 19636 7590 19638 7642
rect 19818 7590 19820 7642
rect 19574 7588 19580 7590
rect 19636 7588 19660 7590
rect 19716 7588 19740 7590
rect 19796 7588 19820 7590
rect 19876 7588 19882 7590
rect 19574 7568 19882 7588
rect 34934 7100 35242 7120
rect 34934 7098 34940 7100
rect 34996 7098 35020 7100
rect 35076 7098 35100 7100
rect 35156 7098 35180 7100
rect 35236 7098 35242 7100
rect 34996 7046 34998 7098
rect 35178 7046 35180 7098
rect 34934 7044 34940 7046
rect 34996 7044 35020 7046
rect 35076 7044 35100 7046
rect 35156 7044 35180 7046
rect 35236 7044 35242 7046
rect 34934 7024 35242 7044
rect 19574 6556 19882 6576
rect 19574 6554 19580 6556
rect 19636 6554 19660 6556
rect 19716 6554 19740 6556
rect 19796 6554 19820 6556
rect 19876 6554 19882 6556
rect 19636 6502 19638 6554
rect 19818 6502 19820 6554
rect 19574 6500 19580 6502
rect 19636 6500 19660 6502
rect 19716 6500 19740 6502
rect 19796 6500 19820 6502
rect 19876 6500 19882 6502
rect 19574 6480 19882 6500
rect 34934 6012 35242 6032
rect 34934 6010 34940 6012
rect 34996 6010 35020 6012
rect 35076 6010 35100 6012
rect 35156 6010 35180 6012
rect 35236 6010 35242 6012
rect 34996 5958 34998 6010
rect 35178 5958 35180 6010
rect 34934 5956 34940 5958
rect 34996 5956 35020 5958
rect 35076 5956 35100 5958
rect 35156 5956 35180 5958
rect 35236 5956 35242 5958
rect 34934 5936 35242 5956
rect 19574 5468 19882 5488
rect 19574 5466 19580 5468
rect 19636 5466 19660 5468
rect 19716 5466 19740 5468
rect 19796 5466 19820 5468
rect 19876 5466 19882 5468
rect 19636 5414 19638 5466
rect 19818 5414 19820 5466
rect 19574 5412 19580 5414
rect 19636 5412 19660 5414
rect 19716 5412 19740 5414
rect 19796 5412 19820 5414
rect 19876 5412 19882 5414
rect 19574 5392 19882 5412
rect 34934 4924 35242 4944
rect 34934 4922 34940 4924
rect 34996 4922 35020 4924
rect 35076 4922 35100 4924
rect 35156 4922 35180 4924
rect 35236 4922 35242 4924
rect 34996 4870 34998 4922
rect 35178 4870 35180 4922
rect 34934 4868 34940 4870
rect 34996 4868 35020 4870
rect 35076 4868 35100 4870
rect 35156 4868 35180 4870
rect 35236 4868 35242 4870
rect 34934 4848 35242 4868
rect 8208 4616 8260 4622
rect 8208 4558 8260 4564
rect 7564 4140 7616 4146
rect 7564 4082 7616 4088
rect 2780 4072 2832 4078
rect 2780 4014 2832 4020
rect 4712 4072 4764 4078
rect 4712 4014 4764 4020
rect 4068 3936 4120 3942
rect 4068 3878 4120 3884
rect 4080 3602 4108 3878
rect 4214 3836 4522 3856
rect 4214 3834 4220 3836
rect 4276 3834 4300 3836
rect 4356 3834 4380 3836
rect 4436 3834 4460 3836
rect 4516 3834 4522 3836
rect 4276 3782 4278 3834
rect 4458 3782 4460 3834
rect 4214 3780 4220 3782
rect 4276 3780 4300 3782
rect 4356 3780 4380 3782
rect 4436 3780 4460 3782
rect 4516 3780 4522 3782
rect 4214 3760 4522 3780
rect 4068 3596 4120 3602
rect 4068 3538 4120 3544
rect 4620 3596 4672 3602
rect 4620 3538 4672 3544
rect 4252 3460 4304 3466
rect 4252 3402 4304 3408
rect 4264 3194 4292 3402
rect 4252 3188 4304 3194
rect 4252 3130 4304 3136
rect 4214 2748 4522 2768
rect 4214 2746 4220 2748
rect 4276 2746 4300 2748
rect 4356 2746 4380 2748
rect 4436 2746 4460 2748
rect 4516 2746 4522 2748
rect 4276 2694 4278 2746
rect 4458 2694 4460 2746
rect 4214 2692 4220 2694
rect 4276 2692 4300 2694
rect 4356 2692 4380 2694
rect 4436 2692 4460 2694
rect 4516 2692 4522 2694
rect 4214 2672 4522 2692
rect 4632 1714 4660 3538
rect 4724 3058 4752 4014
rect 7576 3534 7604 4082
rect 7564 3528 7616 3534
rect 7564 3470 7616 3476
rect 4712 3052 4764 3058
rect 4712 2994 4764 3000
rect 7576 2650 7604 3470
rect 8220 3466 8248 4558
rect 19574 4380 19882 4400
rect 19574 4378 19580 4380
rect 19636 4378 19660 4380
rect 19716 4378 19740 4380
rect 19796 4378 19820 4380
rect 19876 4378 19882 4380
rect 19636 4326 19638 4378
rect 19818 4326 19820 4378
rect 19574 4324 19580 4326
rect 19636 4324 19660 4326
rect 19716 4324 19740 4326
rect 19796 4324 19820 4326
rect 19876 4324 19882 4326
rect 19574 4304 19882 4324
rect 20628 3936 20680 3942
rect 20628 3878 20680 3884
rect 14188 3596 14240 3602
rect 14188 3538 14240 3544
rect 8208 3460 8260 3466
rect 8208 3402 8260 3408
rect 7564 2644 7616 2650
rect 7564 2586 7616 2592
rect 7104 2372 7156 2378
rect 7104 2314 7156 2320
rect 4540 1686 4660 1714
rect 4540 800 4568 1686
rect 7116 800 7144 2314
rect 14200 800 14228 3538
rect 20640 3534 20668 3878
rect 34934 3836 35242 3856
rect 34934 3834 34940 3836
rect 34996 3834 35020 3836
rect 35076 3834 35100 3836
rect 35156 3834 35180 3836
rect 35236 3834 35242 3836
rect 34996 3782 34998 3834
rect 35178 3782 35180 3834
rect 34934 3780 34940 3782
rect 34996 3780 35020 3782
rect 35076 3780 35100 3782
rect 35156 3780 35180 3782
rect 35236 3780 35242 3782
rect 34934 3760 35242 3780
rect 14464 3528 14516 3534
rect 14464 3470 14516 3476
rect 18696 3528 18748 3534
rect 18696 3470 18748 3476
rect 20628 3528 20680 3534
rect 20628 3470 20680 3476
rect 14476 3058 14504 3470
rect 15476 3460 15528 3466
rect 15476 3402 15528 3408
rect 16764 3460 16816 3466
rect 16764 3402 16816 3408
rect 18420 3460 18472 3466
rect 18420 3402 18472 3408
rect 15488 3194 15516 3402
rect 15476 3188 15528 3194
rect 15476 3130 15528 3136
rect 14464 3052 14516 3058
rect 14464 2994 14516 3000
rect 16776 800 16804 3402
rect 18432 3194 18460 3402
rect 18420 3188 18472 3194
rect 18420 3130 18472 3136
rect 18708 3126 18736 3470
rect 20812 3460 20864 3466
rect 20812 3402 20864 3408
rect 21272 3460 21324 3466
rect 21272 3402 21324 3408
rect 19574 3292 19882 3312
rect 19574 3290 19580 3292
rect 19636 3290 19660 3292
rect 19716 3290 19740 3292
rect 19796 3290 19820 3292
rect 19876 3290 19882 3292
rect 19636 3238 19638 3290
rect 19818 3238 19820 3290
rect 19574 3236 19580 3238
rect 19636 3236 19660 3238
rect 19716 3236 19740 3238
rect 19796 3236 19820 3238
rect 19876 3236 19882 3238
rect 19574 3216 19882 3236
rect 20824 3194 20852 3402
rect 20812 3188 20864 3194
rect 20812 3130 20864 3136
rect 18696 3120 18748 3126
rect 18696 3062 18748 3068
rect 19574 2204 19882 2224
rect 19574 2202 19580 2204
rect 19636 2202 19660 2204
rect 19716 2202 19740 2204
rect 19796 2202 19820 2204
rect 19876 2202 19882 2204
rect 19636 2150 19638 2202
rect 19818 2150 19820 2202
rect 19574 2148 19580 2150
rect 19636 2148 19660 2150
rect 19716 2148 19740 2150
rect 19796 2148 19820 2150
rect 19876 2148 19882 2150
rect 19574 2128 19882 2148
rect 21284 800 21312 3402
rect 34934 2748 35242 2768
rect 34934 2746 34940 2748
rect 34996 2746 35020 2748
rect 35076 2746 35100 2748
rect 35156 2746 35180 2748
rect 35236 2746 35242 2748
rect 34996 2694 34998 2746
rect 35178 2694 35180 2746
rect 34934 2692 34940 2694
rect 34996 2692 35020 2694
rect 35076 2692 35100 2694
rect 35156 2692 35180 2694
rect 35236 2692 35242 2694
rect 34934 2672 35242 2692
rect 23848 2440 23900 2446
rect 23848 2382 23900 2388
rect 23860 800 23888 2382
rect 41524 2378 41552 41386
rect 45572 41138 45600 42230
rect 45744 42016 45796 42022
rect 45744 41958 45796 41964
rect 45756 41682 45784 41958
rect 45744 41676 45796 41682
rect 45744 41618 45796 41624
rect 45848 41274 45876 42638
rect 46032 41614 46060 42706
rect 46112 42628 46164 42634
rect 46112 42570 46164 42576
rect 46124 42362 46152 42570
rect 46112 42356 46164 42362
rect 46112 42298 46164 42304
rect 46952 41818 46980 43182
rect 47044 42838 47072 43318
rect 48136 43104 48188 43110
rect 48136 43046 48188 43052
rect 47032 42832 47084 42838
rect 47032 42774 47084 42780
rect 47044 42362 47072 42774
rect 47768 42696 47820 42702
rect 47768 42638 47820 42644
rect 47032 42356 47084 42362
rect 47032 42298 47084 42304
rect 46940 41812 46992 41818
rect 46940 41754 46992 41760
rect 46020 41608 46072 41614
rect 46020 41550 46072 41556
rect 47044 41546 47072 42298
rect 47780 42022 47808 42638
rect 48148 42566 48176 43046
rect 48240 42770 48268 45970
rect 49240 45892 49292 45898
rect 49240 45834 49292 45840
rect 49252 45626 49280 45834
rect 49436 45626 49464 46650
rect 49620 46578 49648 49030
rect 50294 48988 50602 49008
rect 50294 48986 50300 48988
rect 50356 48986 50380 48988
rect 50436 48986 50460 48988
rect 50516 48986 50540 48988
rect 50596 48986 50602 48988
rect 50356 48934 50358 48986
rect 50538 48934 50540 48986
rect 50294 48932 50300 48934
rect 50356 48932 50380 48934
rect 50436 48932 50460 48934
rect 50516 48932 50540 48934
rect 50596 48932 50602 48934
rect 50294 48912 50602 48932
rect 50632 48822 50660 49030
rect 51184 48890 51212 49166
rect 52276 49088 52328 49094
rect 52276 49030 52328 49036
rect 51172 48884 51224 48890
rect 51172 48826 51224 48832
rect 50620 48816 50672 48822
rect 50620 48758 50672 48764
rect 50294 47900 50602 47920
rect 50294 47898 50300 47900
rect 50356 47898 50380 47900
rect 50436 47898 50460 47900
rect 50516 47898 50540 47900
rect 50596 47898 50602 47900
rect 50356 47846 50358 47898
rect 50538 47846 50540 47898
rect 50294 47844 50300 47846
rect 50356 47844 50380 47846
rect 50436 47844 50460 47846
rect 50516 47844 50540 47846
rect 50596 47844 50602 47846
rect 50294 47824 50602 47844
rect 50804 47660 50856 47666
rect 50804 47602 50856 47608
rect 50816 47122 50844 47602
rect 52288 47122 52316 49030
rect 52656 48822 52684 49234
rect 52644 48816 52696 48822
rect 52644 48758 52696 48764
rect 52656 47122 52684 48758
rect 52736 47252 52788 47258
rect 52736 47194 52788 47200
rect 50804 47116 50856 47122
rect 52276 47116 52328 47122
rect 50856 47076 50936 47104
rect 50804 47058 50856 47064
rect 50294 46812 50602 46832
rect 50294 46810 50300 46812
rect 50356 46810 50380 46812
rect 50436 46810 50460 46812
rect 50516 46810 50540 46812
rect 50596 46810 50602 46812
rect 50356 46758 50358 46810
rect 50538 46758 50540 46810
rect 50294 46756 50300 46758
rect 50356 46756 50380 46758
rect 50436 46756 50460 46758
rect 50516 46756 50540 46758
rect 50596 46756 50602 46758
rect 50294 46736 50602 46756
rect 49608 46572 49660 46578
rect 49608 46514 49660 46520
rect 50804 46436 50856 46442
rect 50804 46378 50856 46384
rect 50620 46368 50672 46374
rect 50620 46310 50672 46316
rect 49884 45824 49936 45830
rect 49884 45766 49936 45772
rect 49240 45620 49292 45626
rect 49240 45562 49292 45568
rect 49424 45620 49476 45626
rect 49424 45562 49476 45568
rect 49436 44538 49464 45562
rect 49896 44878 49924 45766
rect 50294 45724 50602 45744
rect 50294 45722 50300 45724
rect 50356 45722 50380 45724
rect 50436 45722 50460 45724
rect 50516 45722 50540 45724
rect 50596 45722 50602 45724
rect 50356 45670 50358 45722
rect 50538 45670 50540 45722
rect 50294 45668 50300 45670
rect 50356 45668 50380 45670
rect 50436 45668 50460 45670
rect 50516 45668 50540 45670
rect 50596 45668 50602 45670
rect 50294 45648 50602 45668
rect 50632 45422 50660 46310
rect 50816 45422 50844 46378
rect 50908 45966 50936 47076
rect 52276 47058 52328 47064
rect 52644 47116 52696 47122
rect 52644 47058 52696 47064
rect 51080 47048 51132 47054
rect 51080 46990 51132 46996
rect 50988 46028 51040 46034
rect 50988 45970 51040 45976
rect 50896 45960 50948 45966
rect 50896 45902 50948 45908
rect 50620 45416 50672 45422
rect 50620 45358 50672 45364
rect 50804 45416 50856 45422
rect 50804 45358 50856 45364
rect 50160 44940 50212 44946
rect 50160 44882 50212 44888
rect 49884 44872 49936 44878
rect 49884 44814 49936 44820
rect 49424 44532 49476 44538
rect 49424 44474 49476 44480
rect 49436 43450 49464 44474
rect 49896 44402 49924 44814
rect 49884 44396 49936 44402
rect 49884 44338 49936 44344
rect 49700 44328 49752 44334
rect 49700 44270 49752 44276
rect 49424 43444 49476 43450
rect 49424 43386 49476 43392
rect 49332 43240 49384 43246
rect 49332 43182 49384 43188
rect 49344 42906 49372 43182
rect 49332 42900 49384 42906
rect 49332 42842 49384 42848
rect 49436 42770 49464 43386
rect 49712 43246 49740 44270
rect 50068 44192 50120 44198
rect 50068 44134 50120 44140
rect 50080 43246 50108 44134
rect 49700 43240 49752 43246
rect 49700 43182 49752 43188
rect 50068 43240 50120 43246
rect 50068 43182 50120 43188
rect 48228 42764 48280 42770
rect 48228 42706 48280 42712
rect 49424 42764 49476 42770
rect 49424 42706 49476 42712
rect 48504 42696 48556 42702
rect 48504 42638 48556 42644
rect 48136 42560 48188 42566
rect 48136 42502 48188 42508
rect 48516 42362 48544 42638
rect 49436 42362 49464 42706
rect 48504 42356 48556 42362
rect 48504 42298 48556 42304
rect 49424 42356 49476 42362
rect 49424 42298 49476 42304
rect 49712 42158 49740 43182
rect 50080 42906 50108 43182
rect 50068 42900 50120 42906
rect 50068 42842 50120 42848
rect 50080 42158 50108 42842
rect 50172 42770 50200 44882
rect 50294 44636 50602 44656
rect 50294 44634 50300 44636
rect 50356 44634 50380 44636
rect 50436 44634 50460 44636
rect 50516 44634 50540 44636
rect 50596 44634 50602 44636
rect 50356 44582 50358 44634
rect 50538 44582 50540 44634
rect 50294 44580 50300 44582
rect 50356 44580 50380 44582
rect 50436 44580 50460 44582
rect 50516 44580 50540 44582
rect 50596 44580 50602 44582
rect 50294 44560 50602 44580
rect 50632 44334 50660 45358
rect 50620 44328 50672 44334
rect 50620 44270 50672 44276
rect 50816 44198 50844 45358
rect 50908 45082 50936 45902
rect 51000 45529 51028 45970
rect 50986 45520 51042 45529
rect 50986 45455 51042 45464
rect 51092 45422 51120 46990
rect 52748 46374 52776 47194
rect 52920 47116 52972 47122
rect 52920 47058 52972 47064
rect 52736 46368 52788 46374
rect 52788 46316 52868 46322
rect 52736 46310 52868 46316
rect 52748 46294 52868 46310
rect 52736 45960 52788 45966
rect 52736 45902 52788 45908
rect 52748 45626 52776 45902
rect 52736 45620 52788 45626
rect 52736 45562 52788 45568
rect 52642 45520 52698 45529
rect 52840 45490 52868 46294
rect 52932 46034 52960 47058
rect 53012 46640 53064 46646
rect 53012 46582 53064 46588
rect 52920 46028 52972 46034
rect 52920 45970 52972 45976
rect 52642 45455 52698 45464
rect 52828 45484 52880 45490
rect 51080 45416 51132 45422
rect 51080 45358 51132 45364
rect 50896 45076 50948 45082
rect 50896 45018 50948 45024
rect 52368 44804 52420 44810
rect 52368 44746 52420 44752
rect 51448 44736 51500 44742
rect 51448 44678 51500 44684
rect 51460 44334 51488 44678
rect 51448 44328 51500 44334
rect 51448 44270 51500 44276
rect 52380 44198 52408 44746
rect 50804 44192 50856 44198
rect 50804 44134 50856 44140
rect 52368 44192 52420 44198
rect 52368 44134 52420 44140
rect 50294 43548 50602 43568
rect 50294 43546 50300 43548
rect 50356 43546 50380 43548
rect 50436 43546 50460 43548
rect 50516 43546 50540 43548
rect 50596 43546 50602 43548
rect 50356 43494 50358 43546
rect 50538 43494 50540 43546
rect 50294 43492 50300 43494
rect 50356 43492 50380 43494
rect 50436 43492 50460 43494
rect 50516 43492 50540 43494
rect 50596 43492 50602 43494
rect 50294 43472 50602 43492
rect 50160 42764 50212 42770
rect 50160 42706 50212 42712
rect 49516 42152 49568 42158
rect 49516 42094 49568 42100
rect 49700 42152 49752 42158
rect 49700 42094 49752 42100
rect 50068 42152 50120 42158
rect 50172 42140 50200 42706
rect 52092 42560 52144 42566
rect 52092 42502 52144 42508
rect 52380 42514 52408 44134
rect 52460 43308 52512 43314
rect 52460 43250 52512 43256
rect 52472 42702 52500 43250
rect 52656 42770 52684 45455
rect 52828 45426 52880 45432
rect 53024 45286 53052 46582
rect 53288 46436 53340 46442
rect 53288 46378 53340 46384
rect 53300 46102 53328 46378
rect 53288 46096 53340 46102
rect 53288 46038 53340 46044
rect 53196 46028 53248 46034
rect 53196 45970 53248 45976
rect 53208 45529 53236 45970
rect 53300 45626 53328 46038
rect 53288 45620 53340 45626
rect 53288 45562 53340 45568
rect 53194 45520 53250 45529
rect 53194 45455 53250 45464
rect 53012 45280 53064 45286
rect 53012 45222 53064 45228
rect 52736 44736 52788 44742
rect 52736 44678 52788 44684
rect 52748 44470 52776 44678
rect 53024 44538 53052 45222
rect 53012 44532 53064 44538
rect 53012 44474 53064 44480
rect 52736 44464 52788 44470
rect 52736 44406 52788 44412
rect 53012 44396 53064 44402
rect 53012 44338 53064 44344
rect 53024 43450 53052 44338
rect 53012 43444 53064 43450
rect 53012 43386 53064 43392
rect 52828 43308 52880 43314
rect 52828 43250 52880 43256
rect 52736 43104 52788 43110
rect 52736 43046 52788 43052
rect 52644 42764 52696 42770
rect 52644 42706 52696 42712
rect 52460 42696 52512 42702
rect 52460 42638 52512 42644
rect 52552 42696 52604 42702
rect 52552 42638 52604 42644
rect 52564 42514 52592 42638
rect 50294 42460 50602 42480
rect 50294 42458 50300 42460
rect 50356 42458 50380 42460
rect 50436 42458 50460 42460
rect 50516 42458 50540 42460
rect 50596 42458 50602 42460
rect 50356 42406 50358 42458
rect 50538 42406 50540 42458
rect 50294 42404 50300 42406
rect 50356 42404 50380 42406
rect 50436 42404 50460 42406
rect 50516 42404 50540 42406
rect 50596 42404 50602 42406
rect 50294 42384 50602 42404
rect 52000 42356 52052 42362
rect 52104 42344 52132 42502
rect 52380 42486 52592 42514
rect 52052 42316 52132 42344
rect 52000 42298 52052 42304
rect 50344 42152 50396 42158
rect 50172 42112 50344 42140
rect 50068 42094 50120 42100
rect 50344 42094 50396 42100
rect 51080 42152 51132 42158
rect 51080 42094 51132 42100
rect 51724 42152 51776 42158
rect 51724 42094 51776 42100
rect 47768 42016 47820 42022
rect 47768 41958 47820 41964
rect 47124 41812 47176 41818
rect 47124 41754 47176 41760
rect 47032 41540 47084 41546
rect 47032 41482 47084 41488
rect 45836 41268 45888 41274
rect 45836 41210 45888 41216
rect 47136 41138 47164 41754
rect 49528 41546 49556 42094
rect 50080 42022 50108 42094
rect 50068 42016 50120 42022
rect 50068 41958 50120 41964
rect 51092 41682 51120 42094
rect 51736 41682 51764 42094
rect 52748 41818 52776 43046
rect 52840 42362 52868 43250
rect 52920 43240 52972 43246
rect 52920 43182 52972 43188
rect 52932 42362 52960 43182
rect 53012 43172 53064 43178
rect 53012 43114 53064 43120
rect 52828 42356 52880 42362
rect 52828 42298 52880 42304
rect 52920 42356 52972 42362
rect 52920 42298 52972 42304
rect 53024 42226 53052 43114
rect 53656 42560 53708 42566
rect 53656 42502 53708 42508
rect 53012 42220 53064 42226
rect 53012 42162 53064 42168
rect 52736 41812 52788 41818
rect 52736 41754 52788 41760
rect 51080 41676 51132 41682
rect 51080 41618 51132 41624
rect 51724 41676 51776 41682
rect 51724 41618 51776 41624
rect 53668 41614 53696 42502
rect 53656 41608 53708 41614
rect 53656 41550 53708 41556
rect 49516 41540 49568 41546
rect 49516 41482 49568 41488
rect 50294 41372 50602 41392
rect 50294 41370 50300 41372
rect 50356 41370 50380 41372
rect 50436 41370 50460 41372
rect 50516 41370 50540 41372
rect 50596 41370 50602 41372
rect 50356 41318 50358 41370
rect 50538 41318 50540 41370
rect 50294 41316 50300 41318
rect 50356 41316 50380 41318
rect 50436 41316 50460 41318
rect 50516 41316 50540 41318
rect 50596 41316 50602 41318
rect 50294 41296 50602 41316
rect 45560 41132 45612 41138
rect 45560 41074 45612 41080
rect 47124 41132 47176 41138
rect 47124 41074 47176 41080
rect 50294 40284 50602 40304
rect 50294 40282 50300 40284
rect 50356 40282 50380 40284
rect 50436 40282 50460 40284
rect 50516 40282 50540 40284
rect 50596 40282 50602 40284
rect 50356 40230 50358 40282
rect 50538 40230 50540 40282
rect 50294 40228 50300 40230
rect 50356 40228 50380 40230
rect 50436 40228 50460 40230
rect 50516 40228 50540 40230
rect 50596 40228 50602 40230
rect 50294 40208 50602 40228
rect 50294 39196 50602 39216
rect 50294 39194 50300 39196
rect 50356 39194 50380 39196
rect 50436 39194 50460 39196
rect 50516 39194 50540 39196
rect 50596 39194 50602 39196
rect 50356 39142 50358 39194
rect 50538 39142 50540 39194
rect 50294 39140 50300 39142
rect 50356 39140 50380 39142
rect 50436 39140 50460 39142
rect 50516 39140 50540 39142
rect 50596 39140 50602 39142
rect 50294 39120 50602 39140
rect 50294 38108 50602 38128
rect 50294 38106 50300 38108
rect 50356 38106 50380 38108
rect 50436 38106 50460 38108
rect 50516 38106 50540 38108
rect 50596 38106 50602 38108
rect 50356 38054 50358 38106
rect 50538 38054 50540 38106
rect 50294 38052 50300 38054
rect 50356 38052 50380 38054
rect 50436 38052 50460 38054
rect 50516 38052 50540 38054
rect 50596 38052 50602 38054
rect 50294 38032 50602 38052
rect 50294 37020 50602 37040
rect 50294 37018 50300 37020
rect 50356 37018 50380 37020
rect 50436 37018 50460 37020
rect 50516 37018 50540 37020
rect 50596 37018 50602 37020
rect 50356 36966 50358 37018
rect 50538 36966 50540 37018
rect 50294 36964 50300 36966
rect 50356 36964 50380 36966
rect 50436 36964 50460 36966
rect 50516 36964 50540 36966
rect 50596 36964 50602 36966
rect 50294 36944 50602 36964
rect 50294 35932 50602 35952
rect 50294 35930 50300 35932
rect 50356 35930 50380 35932
rect 50436 35930 50460 35932
rect 50516 35930 50540 35932
rect 50596 35930 50602 35932
rect 50356 35878 50358 35930
rect 50538 35878 50540 35930
rect 50294 35876 50300 35878
rect 50356 35876 50380 35878
rect 50436 35876 50460 35878
rect 50516 35876 50540 35878
rect 50596 35876 50602 35878
rect 50294 35856 50602 35876
rect 55600 35894 55628 55626
rect 56232 55412 56284 55418
rect 56232 55354 56284 55360
rect 55600 35866 55720 35894
rect 50294 34844 50602 34864
rect 50294 34842 50300 34844
rect 50356 34842 50380 34844
rect 50436 34842 50460 34844
rect 50516 34842 50540 34844
rect 50596 34842 50602 34844
rect 50356 34790 50358 34842
rect 50538 34790 50540 34842
rect 50294 34788 50300 34790
rect 50356 34788 50380 34790
rect 50436 34788 50460 34790
rect 50516 34788 50540 34790
rect 50596 34788 50602 34790
rect 50294 34768 50602 34788
rect 50294 33756 50602 33776
rect 50294 33754 50300 33756
rect 50356 33754 50380 33756
rect 50436 33754 50460 33756
rect 50516 33754 50540 33756
rect 50596 33754 50602 33756
rect 50356 33702 50358 33754
rect 50538 33702 50540 33754
rect 50294 33700 50300 33702
rect 50356 33700 50380 33702
rect 50436 33700 50460 33702
rect 50516 33700 50540 33702
rect 50596 33700 50602 33702
rect 50294 33680 50602 33700
rect 50294 32668 50602 32688
rect 50294 32666 50300 32668
rect 50356 32666 50380 32668
rect 50436 32666 50460 32668
rect 50516 32666 50540 32668
rect 50596 32666 50602 32668
rect 50356 32614 50358 32666
rect 50538 32614 50540 32666
rect 50294 32612 50300 32614
rect 50356 32612 50380 32614
rect 50436 32612 50460 32614
rect 50516 32612 50540 32614
rect 50596 32612 50602 32614
rect 50294 32592 50602 32612
rect 50294 31580 50602 31600
rect 50294 31578 50300 31580
rect 50356 31578 50380 31580
rect 50436 31578 50460 31580
rect 50516 31578 50540 31580
rect 50596 31578 50602 31580
rect 50356 31526 50358 31578
rect 50538 31526 50540 31578
rect 50294 31524 50300 31526
rect 50356 31524 50380 31526
rect 50436 31524 50460 31526
rect 50516 31524 50540 31526
rect 50596 31524 50602 31526
rect 50294 31504 50602 31524
rect 50294 30492 50602 30512
rect 50294 30490 50300 30492
rect 50356 30490 50380 30492
rect 50436 30490 50460 30492
rect 50516 30490 50540 30492
rect 50596 30490 50602 30492
rect 50356 30438 50358 30490
rect 50538 30438 50540 30490
rect 50294 30436 50300 30438
rect 50356 30436 50380 30438
rect 50436 30436 50460 30438
rect 50516 30436 50540 30438
rect 50596 30436 50602 30438
rect 50294 30416 50602 30436
rect 50294 29404 50602 29424
rect 50294 29402 50300 29404
rect 50356 29402 50380 29404
rect 50436 29402 50460 29404
rect 50516 29402 50540 29404
rect 50596 29402 50602 29404
rect 50356 29350 50358 29402
rect 50538 29350 50540 29402
rect 50294 29348 50300 29350
rect 50356 29348 50380 29350
rect 50436 29348 50460 29350
rect 50516 29348 50540 29350
rect 50596 29348 50602 29350
rect 50294 29328 50602 29348
rect 50294 28316 50602 28336
rect 50294 28314 50300 28316
rect 50356 28314 50380 28316
rect 50436 28314 50460 28316
rect 50516 28314 50540 28316
rect 50596 28314 50602 28316
rect 50356 28262 50358 28314
rect 50538 28262 50540 28314
rect 50294 28260 50300 28262
rect 50356 28260 50380 28262
rect 50436 28260 50460 28262
rect 50516 28260 50540 28262
rect 50596 28260 50602 28262
rect 50294 28240 50602 28260
rect 50294 27228 50602 27248
rect 50294 27226 50300 27228
rect 50356 27226 50380 27228
rect 50436 27226 50460 27228
rect 50516 27226 50540 27228
rect 50596 27226 50602 27228
rect 50356 27174 50358 27226
rect 50538 27174 50540 27226
rect 50294 27172 50300 27174
rect 50356 27172 50380 27174
rect 50436 27172 50460 27174
rect 50516 27172 50540 27174
rect 50596 27172 50602 27174
rect 50294 27152 50602 27172
rect 50294 26140 50602 26160
rect 50294 26138 50300 26140
rect 50356 26138 50380 26140
rect 50436 26138 50460 26140
rect 50516 26138 50540 26140
rect 50596 26138 50602 26140
rect 50356 26086 50358 26138
rect 50538 26086 50540 26138
rect 50294 26084 50300 26086
rect 50356 26084 50380 26086
rect 50436 26084 50460 26086
rect 50516 26084 50540 26086
rect 50596 26084 50602 26086
rect 50294 26064 50602 26084
rect 50294 25052 50602 25072
rect 50294 25050 50300 25052
rect 50356 25050 50380 25052
rect 50436 25050 50460 25052
rect 50516 25050 50540 25052
rect 50596 25050 50602 25052
rect 50356 24998 50358 25050
rect 50538 24998 50540 25050
rect 50294 24996 50300 24998
rect 50356 24996 50380 24998
rect 50436 24996 50460 24998
rect 50516 24996 50540 24998
rect 50596 24996 50602 24998
rect 50294 24976 50602 24996
rect 50294 23964 50602 23984
rect 50294 23962 50300 23964
rect 50356 23962 50380 23964
rect 50436 23962 50460 23964
rect 50516 23962 50540 23964
rect 50596 23962 50602 23964
rect 50356 23910 50358 23962
rect 50538 23910 50540 23962
rect 50294 23908 50300 23910
rect 50356 23908 50380 23910
rect 50436 23908 50460 23910
rect 50516 23908 50540 23910
rect 50596 23908 50602 23910
rect 50294 23888 50602 23908
rect 55692 23526 55720 35866
rect 56244 24750 56272 55354
rect 56324 42696 56376 42702
rect 56324 42638 56376 42644
rect 56336 41682 56364 42638
rect 56888 42226 56916 55694
rect 58164 47048 58216 47054
rect 58162 47016 58164 47025
rect 58216 47016 58218 47025
rect 58162 46951 58218 46960
rect 57060 42628 57112 42634
rect 57060 42570 57112 42576
rect 56876 42220 56928 42226
rect 56876 42162 56928 42168
rect 56508 42016 56560 42022
rect 56508 41958 56560 41964
rect 56520 41682 56548 41958
rect 56324 41676 56376 41682
rect 56324 41618 56376 41624
rect 56508 41676 56560 41682
rect 56508 41618 56560 41624
rect 57072 31890 57100 42570
rect 58162 42256 58218 42265
rect 58162 42191 58218 42200
rect 58176 41682 58204 42191
rect 58164 41676 58216 41682
rect 58164 41618 58216 41624
rect 58162 32056 58218 32065
rect 58162 31991 58218 32000
rect 57060 31884 57112 31890
rect 57060 31826 57112 31832
rect 58176 31822 58204 31991
rect 58164 31816 58216 31822
rect 58164 31758 58216 31764
rect 57702 29336 57758 29345
rect 57702 29271 57758 29280
rect 56968 29164 57020 29170
rect 56968 29106 57020 29112
rect 56232 24744 56284 24750
rect 56232 24686 56284 24692
rect 55680 23520 55732 23526
rect 55680 23462 55732 23468
rect 50294 22876 50602 22896
rect 50294 22874 50300 22876
rect 50356 22874 50380 22876
rect 50436 22874 50460 22876
rect 50516 22874 50540 22876
rect 50596 22874 50602 22876
rect 50356 22822 50358 22874
rect 50538 22822 50540 22874
rect 50294 22820 50300 22822
rect 50356 22820 50380 22822
rect 50436 22820 50460 22822
rect 50516 22820 50540 22822
rect 50596 22820 50602 22822
rect 50294 22800 50602 22820
rect 50294 21788 50602 21808
rect 50294 21786 50300 21788
rect 50356 21786 50380 21788
rect 50436 21786 50460 21788
rect 50516 21786 50540 21788
rect 50596 21786 50602 21788
rect 50356 21734 50358 21786
rect 50538 21734 50540 21786
rect 50294 21732 50300 21734
rect 50356 21732 50380 21734
rect 50436 21732 50460 21734
rect 50516 21732 50540 21734
rect 50596 21732 50602 21734
rect 50294 21712 50602 21732
rect 50294 20700 50602 20720
rect 50294 20698 50300 20700
rect 50356 20698 50380 20700
rect 50436 20698 50460 20700
rect 50516 20698 50540 20700
rect 50596 20698 50602 20700
rect 50356 20646 50358 20698
rect 50538 20646 50540 20698
rect 50294 20644 50300 20646
rect 50356 20644 50380 20646
rect 50436 20644 50460 20646
rect 50516 20644 50540 20646
rect 50596 20644 50602 20646
rect 50294 20624 50602 20644
rect 50294 19612 50602 19632
rect 50294 19610 50300 19612
rect 50356 19610 50380 19612
rect 50436 19610 50460 19612
rect 50516 19610 50540 19612
rect 50596 19610 50602 19612
rect 50356 19558 50358 19610
rect 50538 19558 50540 19610
rect 50294 19556 50300 19558
rect 50356 19556 50380 19558
rect 50436 19556 50460 19558
rect 50516 19556 50540 19558
rect 50596 19556 50602 19558
rect 50294 19536 50602 19556
rect 50294 18524 50602 18544
rect 50294 18522 50300 18524
rect 50356 18522 50380 18524
rect 50436 18522 50460 18524
rect 50516 18522 50540 18524
rect 50596 18522 50602 18524
rect 50356 18470 50358 18522
rect 50538 18470 50540 18522
rect 50294 18468 50300 18470
rect 50356 18468 50380 18470
rect 50436 18468 50460 18470
rect 50516 18468 50540 18470
rect 50596 18468 50602 18470
rect 50294 18448 50602 18468
rect 50294 17436 50602 17456
rect 50294 17434 50300 17436
rect 50356 17434 50380 17436
rect 50436 17434 50460 17436
rect 50516 17434 50540 17436
rect 50596 17434 50602 17436
rect 50356 17382 50358 17434
rect 50538 17382 50540 17434
rect 50294 17380 50300 17382
rect 50356 17380 50380 17382
rect 50436 17380 50460 17382
rect 50516 17380 50540 17382
rect 50596 17380 50602 17382
rect 50294 17360 50602 17380
rect 50294 16348 50602 16368
rect 50294 16346 50300 16348
rect 50356 16346 50380 16348
rect 50436 16346 50460 16348
rect 50516 16346 50540 16348
rect 50596 16346 50602 16348
rect 50356 16294 50358 16346
rect 50538 16294 50540 16346
rect 50294 16292 50300 16294
rect 50356 16292 50380 16294
rect 50436 16292 50460 16294
rect 50516 16292 50540 16294
rect 50596 16292 50602 16294
rect 50294 16272 50602 16292
rect 50294 15260 50602 15280
rect 50294 15258 50300 15260
rect 50356 15258 50380 15260
rect 50436 15258 50460 15260
rect 50516 15258 50540 15260
rect 50596 15258 50602 15260
rect 50356 15206 50358 15258
rect 50538 15206 50540 15258
rect 50294 15204 50300 15206
rect 50356 15204 50380 15206
rect 50436 15204 50460 15206
rect 50516 15204 50540 15206
rect 50596 15204 50602 15206
rect 50294 15184 50602 15204
rect 50294 14172 50602 14192
rect 50294 14170 50300 14172
rect 50356 14170 50380 14172
rect 50436 14170 50460 14172
rect 50516 14170 50540 14172
rect 50596 14170 50602 14172
rect 50356 14118 50358 14170
rect 50538 14118 50540 14170
rect 50294 14116 50300 14118
rect 50356 14116 50380 14118
rect 50436 14116 50460 14118
rect 50516 14116 50540 14118
rect 50596 14116 50602 14118
rect 50294 14096 50602 14116
rect 50294 13084 50602 13104
rect 50294 13082 50300 13084
rect 50356 13082 50380 13084
rect 50436 13082 50460 13084
rect 50516 13082 50540 13084
rect 50596 13082 50602 13084
rect 50356 13030 50358 13082
rect 50538 13030 50540 13082
rect 50294 13028 50300 13030
rect 50356 13028 50380 13030
rect 50436 13028 50460 13030
rect 50516 13028 50540 13030
rect 50596 13028 50602 13030
rect 50294 13008 50602 13028
rect 50294 11996 50602 12016
rect 50294 11994 50300 11996
rect 50356 11994 50380 11996
rect 50436 11994 50460 11996
rect 50516 11994 50540 11996
rect 50596 11994 50602 11996
rect 50356 11942 50358 11994
rect 50538 11942 50540 11994
rect 50294 11940 50300 11942
rect 50356 11940 50380 11942
rect 50436 11940 50460 11942
rect 50516 11940 50540 11942
rect 50596 11940 50602 11942
rect 50294 11920 50602 11940
rect 50294 10908 50602 10928
rect 50294 10906 50300 10908
rect 50356 10906 50380 10908
rect 50436 10906 50460 10908
rect 50516 10906 50540 10908
rect 50596 10906 50602 10908
rect 50356 10854 50358 10906
rect 50538 10854 50540 10906
rect 50294 10852 50300 10854
rect 50356 10852 50380 10854
rect 50436 10852 50460 10854
rect 50516 10852 50540 10854
rect 50596 10852 50602 10854
rect 50294 10832 50602 10852
rect 50294 9820 50602 9840
rect 50294 9818 50300 9820
rect 50356 9818 50380 9820
rect 50436 9818 50460 9820
rect 50516 9818 50540 9820
rect 50596 9818 50602 9820
rect 50356 9766 50358 9818
rect 50538 9766 50540 9818
rect 50294 9764 50300 9766
rect 50356 9764 50380 9766
rect 50436 9764 50460 9766
rect 50516 9764 50540 9766
rect 50596 9764 50602 9766
rect 50294 9744 50602 9764
rect 50294 8732 50602 8752
rect 50294 8730 50300 8732
rect 50356 8730 50380 8732
rect 50436 8730 50460 8732
rect 50516 8730 50540 8732
rect 50596 8730 50602 8732
rect 50356 8678 50358 8730
rect 50538 8678 50540 8730
rect 50294 8676 50300 8678
rect 50356 8676 50380 8678
rect 50436 8676 50460 8678
rect 50516 8676 50540 8678
rect 50596 8676 50602 8678
rect 50294 8656 50602 8676
rect 50294 7644 50602 7664
rect 50294 7642 50300 7644
rect 50356 7642 50380 7644
rect 50436 7642 50460 7644
rect 50516 7642 50540 7644
rect 50596 7642 50602 7644
rect 50356 7590 50358 7642
rect 50538 7590 50540 7642
rect 50294 7588 50300 7590
rect 50356 7588 50380 7590
rect 50436 7588 50460 7590
rect 50516 7588 50540 7590
rect 50596 7588 50602 7590
rect 50294 7568 50602 7588
rect 50294 6556 50602 6576
rect 50294 6554 50300 6556
rect 50356 6554 50380 6556
rect 50436 6554 50460 6556
rect 50516 6554 50540 6556
rect 50596 6554 50602 6556
rect 50356 6502 50358 6554
rect 50538 6502 50540 6554
rect 50294 6500 50300 6502
rect 50356 6500 50380 6502
rect 50436 6500 50460 6502
rect 50516 6500 50540 6502
rect 50596 6500 50602 6502
rect 50294 6480 50602 6500
rect 50294 5468 50602 5488
rect 50294 5466 50300 5468
rect 50356 5466 50380 5468
rect 50436 5466 50460 5468
rect 50516 5466 50540 5468
rect 50596 5466 50602 5468
rect 50356 5414 50358 5466
rect 50538 5414 50540 5466
rect 50294 5412 50300 5414
rect 50356 5412 50380 5414
rect 50436 5412 50460 5414
rect 50516 5412 50540 5414
rect 50596 5412 50602 5414
rect 50294 5392 50602 5412
rect 50294 4380 50602 4400
rect 50294 4378 50300 4380
rect 50356 4378 50380 4380
rect 50436 4378 50460 4380
rect 50516 4378 50540 4380
rect 50596 4378 50602 4380
rect 50356 4326 50358 4378
rect 50538 4326 50540 4378
rect 50294 4324 50300 4326
rect 50356 4324 50380 4326
rect 50436 4324 50460 4326
rect 50516 4324 50540 4326
rect 50596 4324 50602 4326
rect 50294 4304 50602 4324
rect 51448 4072 51500 4078
rect 51448 4014 51500 4020
rect 45192 3596 45244 3602
rect 45192 3538 45244 3544
rect 44640 3528 44692 3534
rect 45204 3482 45232 3538
rect 44640 3470 44692 3476
rect 44652 3058 44680 3470
rect 45112 3454 45232 3482
rect 44640 3052 44692 3058
rect 44640 2994 44692 3000
rect 41512 2372 41564 2378
rect 41512 2314 41564 2320
rect 45112 800 45140 3454
rect 50160 3392 50212 3398
rect 50160 3334 50212 3340
rect 50172 2922 50200 3334
rect 50294 3292 50602 3312
rect 50294 3290 50300 3292
rect 50356 3290 50380 3292
rect 50436 3290 50460 3292
rect 50516 3290 50540 3292
rect 50596 3290 50602 3292
rect 50356 3238 50358 3290
rect 50538 3238 50540 3290
rect 50294 3236 50300 3238
rect 50356 3236 50380 3238
rect 50436 3236 50460 3238
rect 50516 3236 50540 3238
rect 50596 3236 50602 3238
rect 50294 3216 50602 3236
rect 51460 3058 51488 4014
rect 51540 3936 51592 3942
rect 51540 3878 51592 3884
rect 54484 3936 54536 3942
rect 54484 3878 54536 3884
rect 51552 3602 51580 3878
rect 51540 3596 51592 3602
rect 51540 3538 51592 3544
rect 52184 3596 52236 3602
rect 52184 3538 52236 3544
rect 51724 3460 51776 3466
rect 51724 3402 51776 3408
rect 51736 3194 51764 3402
rect 51724 3188 51776 3194
rect 51724 3130 51776 3136
rect 51448 3052 51500 3058
rect 51448 2994 51500 3000
rect 50160 2916 50212 2922
rect 50160 2858 50212 2864
rect 50294 2204 50602 2224
rect 50294 2202 50300 2204
rect 50356 2202 50380 2204
rect 50436 2202 50460 2204
rect 50516 2202 50540 2204
rect 50596 2202 50602 2204
rect 50356 2150 50358 2202
rect 50538 2150 50540 2202
rect 50294 2148 50300 2150
rect 50356 2148 50380 2150
rect 50436 2148 50460 2150
rect 50516 2148 50540 2150
rect 50596 2148 50602 2150
rect 50294 2128 50602 2148
rect 52196 800 52224 3538
rect 54496 3058 54524 3878
rect 55692 3534 55720 23462
rect 56140 19372 56192 19378
rect 56140 19314 56192 19320
rect 55680 3528 55732 3534
rect 55680 3470 55732 3476
rect 54668 3392 54720 3398
rect 54668 3334 54720 3340
rect 54680 3126 54708 3334
rect 56152 3194 56180 19314
rect 56244 8498 56272 24686
rect 56508 24608 56560 24614
rect 56508 24550 56560 24556
rect 56520 24274 56548 24550
rect 56508 24268 56560 24274
rect 56508 24210 56560 24216
rect 56980 22438 57008 29106
rect 57716 28626 57744 29271
rect 57980 29028 58032 29034
rect 57980 28970 58032 28976
rect 57992 28626 58020 28970
rect 58164 28960 58216 28966
rect 58164 28902 58216 28908
rect 58176 28626 58204 28902
rect 57704 28620 57756 28626
rect 57704 28562 57756 28568
rect 57980 28620 58032 28626
rect 57980 28562 58032 28568
rect 58164 28620 58216 28626
rect 58164 28562 58216 28568
rect 57060 24812 57112 24818
rect 57060 24754 57112 24760
rect 57072 23798 57100 24754
rect 57796 24676 57848 24682
rect 57796 24618 57848 24624
rect 57060 23792 57112 23798
rect 57060 23734 57112 23740
rect 56968 22432 57020 22438
rect 56968 22374 57020 22380
rect 56508 19168 56560 19174
rect 56508 19110 56560 19116
rect 56520 18834 56548 19110
rect 56508 18828 56560 18834
rect 56508 18770 56560 18776
rect 56324 12232 56376 12238
rect 56324 12174 56376 12180
rect 56336 11218 56364 12174
rect 56980 11762 57008 22374
rect 56968 11756 57020 11762
rect 56968 11698 57020 11704
rect 56508 11552 56560 11558
rect 56508 11494 56560 11500
rect 56520 11218 56548 11494
rect 56324 11212 56376 11218
rect 56324 11154 56376 11160
rect 56508 11212 56560 11218
rect 56508 11154 56560 11160
rect 56508 8900 56560 8906
rect 56508 8842 56560 8848
rect 56520 8634 56548 8842
rect 56508 8628 56560 8634
rect 56508 8570 56560 8576
rect 56232 8492 56284 8498
rect 56232 8434 56284 8440
rect 56140 3188 56192 3194
rect 56140 3130 56192 3136
rect 54668 3120 54720 3126
rect 54668 3062 54720 3068
rect 54484 3052 54536 3058
rect 54484 2994 54536 3000
rect 54760 2984 54812 2990
rect 54760 2926 54812 2932
rect 54772 800 54800 2926
rect 56244 2922 56272 8434
rect 56324 4616 56376 4622
rect 56324 4558 56376 4564
rect 56336 3618 56364 4558
rect 56508 4548 56560 4554
rect 56508 4490 56560 4496
rect 56520 3738 56548 4490
rect 57808 4146 57836 24618
rect 57888 24608 57940 24614
rect 57888 24550 57940 24556
rect 58162 24576 58218 24585
rect 57900 24342 57928 24550
rect 58162 24511 58218 24520
rect 57888 24336 57940 24342
rect 57888 24278 57940 24284
rect 58176 24274 58204 24511
rect 58164 24268 58216 24274
rect 58164 24210 58216 24216
rect 57888 19168 57940 19174
rect 57888 19110 57940 19116
rect 58162 19136 58218 19145
rect 57900 18902 57928 19110
rect 58162 19071 58218 19080
rect 57888 18896 57940 18902
rect 57888 18838 57940 18844
rect 58176 18834 58204 19071
rect 58164 18828 58216 18834
rect 58164 18770 58216 18776
rect 58162 11656 58218 11665
rect 58162 11591 58218 11600
rect 58176 11218 58204 11591
rect 58164 11212 58216 11218
rect 58164 11154 58216 11160
rect 57888 9036 57940 9042
rect 57888 8978 57940 8984
rect 57900 8498 57928 8978
rect 58162 8936 58218 8945
rect 58162 8871 58164 8880
rect 58216 8871 58218 8880
rect 58164 8842 58216 8848
rect 57888 8492 57940 8498
rect 57888 8434 57940 8440
rect 59268 4548 59320 4554
rect 59268 4490 59320 4496
rect 57796 4140 57848 4146
rect 57796 4082 57848 4088
rect 57336 4072 57388 4078
rect 57336 4014 57388 4020
rect 57244 3936 57296 3942
rect 57244 3878 57296 3884
rect 56508 3732 56560 3738
rect 56508 3674 56560 3680
rect 56784 3664 56836 3670
rect 56336 3590 56456 3618
rect 56784 3606 56836 3612
rect 56324 3528 56376 3534
rect 56324 3470 56376 3476
rect 56336 3126 56364 3470
rect 56324 3120 56376 3126
rect 56324 3062 56376 3068
rect 56232 2916 56284 2922
rect 56232 2858 56284 2864
rect 56428 2582 56456 3590
rect 56796 3058 56824 3606
rect 56876 3460 56928 3466
rect 56876 3402 56928 3408
rect 56888 3194 56916 3402
rect 56876 3188 56928 3194
rect 56876 3130 56928 3136
rect 56784 3052 56836 3058
rect 56784 2994 56836 3000
rect 56416 2576 56468 2582
rect 56416 2518 56468 2524
rect 57256 2122 57284 3878
rect 57348 2650 57376 4014
rect 57888 3596 57940 3602
rect 57888 3538 57940 3544
rect 57336 2644 57388 2650
rect 57336 2586 57388 2592
rect 57256 2094 57376 2122
rect 57348 800 57376 2094
rect 57900 1465 57928 3538
rect 57886 1456 57942 1465
rect 57886 1391 57942 1400
rect 59280 800 59308 4490
rect -10 0 102 800
rect 1922 0 2034 800
rect 4498 0 4610 800
rect 7074 0 7186 800
rect 9006 0 9118 800
rect 11582 0 11694 800
rect 14158 0 14270 800
rect 16734 0 16846 800
rect 18666 0 18778 800
rect 21242 0 21354 800
rect 23818 0 23930 800
rect 25750 0 25862 800
rect 28326 0 28438 800
rect 30902 0 31014 800
rect 33478 0 33590 800
rect 35410 0 35522 800
rect 37986 0 38098 800
rect 40562 0 40674 800
rect 42494 0 42606 800
rect 45070 0 45182 800
rect 47646 0 47758 800
rect 50222 0 50334 800
rect 52154 0 52266 800
rect 54730 0 54842 800
rect 57306 0 57418 800
rect 59238 0 59350 800
<< via2 >>
rect 4220 57146 4276 57148
rect 4300 57146 4356 57148
rect 4380 57146 4436 57148
rect 4460 57146 4516 57148
rect 4220 57094 4266 57146
rect 4266 57094 4276 57146
rect 4300 57094 4330 57146
rect 4330 57094 4342 57146
rect 4342 57094 4356 57146
rect 4380 57094 4394 57146
rect 4394 57094 4406 57146
rect 4406 57094 4436 57146
rect 4460 57094 4470 57146
rect 4470 57094 4516 57146
rect 4220 57092 4276 57094
rect 4300 57092 4356 57094
rect 4380 57092 4436 57094
rect 4460 57092 4516 57094
rect 19580 57690 19636 57692
rect 19660 57690 19716 57692
rect 19740 57690 19796 57692
rect 19820 57690 19876 57692
rect 19580 57638 19626 57690
rect 19626 57638 19636 57690
rect 19660 57638 19690 57690
rect 19690 57638 19702 57690
rect 19702 57638 19716 57690
rect 19740 57638 19754 57690
rect 19754 57638 19766 57690
rect 19766 57638 19796 57690
rect 19820 57638 19830 57690
rect 19830 57638 19876 57690
rect 19580 57636 19636 57638
rect 19660 57636 19716 57638
rect 19740 57636 19796 57638
rect 19820 57636 19876 57638
rect 19580 56602 19636 56604
rect 19660 56602 19716 56604
rect 19740 56602 19796 56604
rect 19820 56602 19876 56604
rect 19580 56550 19626 56602
rect 19626 56550 19636 56602
rect 19660 56550 19690 56602
rect 19690 56550 19702 56602
rect 19702 56550 19716 56602
rect 19740 56550 19754 56602
rect 19754 56550 19766 56602
rect 19766 56550 19796 56602
rect 19820 56550 19830 56602
rect 19830 56550 19876 56602
rect 19580 56548 19636 56550
rect 19660 56548 19716 56550
rect 19740 56548 19796 56550
rect 19820 56548 19876 56550
rect 4220 56058 4276 56060
rect 4300 56058 4356 56060
rect 4380 56058 4436 56060
rect 4460 56058 4516 56060
rect 4220 56006 4266 56058
rect 4266 56006 4276 56058
rect 4300 56006 4330 56058
rect 4330 56006 4342 56058
rect 4342 56006 4356 56058
rect 4380 56006 4394 56058
rect 4394 56006 4406 56058
rect 4406 56006 4436 56058
rect 4460 56006 4470 56058
rect 4470 56006 4516 56058
rect 4220 56004 4276 56006
rect 4300 56004 4356 56006
rect 4380 56004 4436 56006
rect 4460 56004 4516 56006
rect 2778 55120 2834 55176
rect 4220 54970 4276 54972
rect 4300 54970 4356 54972
rect 4380 54970 4436 54972
rect 4460 54970 4516 54972
rect 4220 54918 4266 54970
rect 4266 54918 4276 54970
rect 4300 54918 4330 54970
rect 4330 54918 4342 54970
rect 4342 54918 4356 54970
rect 4380 54918 4394 54970
rect 4394 54918 4406 54970
rect 4406 54918 4436 54970
rect 4460 54918 4470 54970
rect 4470 54918 4516 54970
rect 4220 54916 4276 54918
rect 4300 54916 4356 54918
rect 4380 54916 4436 54918
rect 4460 54916 4516 54918
rect 4220 53882 4276 53884
rect 4300 53882 4356 53884
rect 4380 53882 4436 53884
rect 4460 53882 4516 53884
rect 4220 53830 4266 53882
rect 4266 53830 4276 53882
rect 4300 53830 4330 53882
rect 4330 53830 4342 53882
rect 4342 53830 4356 53882
rect 4380 53830 4394 53882
rect 4394 53830 4406 53882
rect 4406 53830 4436 53882
rect 4460 53830 4470 53882
rect 4470 53830 4516 53882
rect 4220 53828 4276 53830
rect 4300 53828 4356 53830
rect 4380 53828 4436 53830
rect 4460 53828 4516 53830
rect 4220 52794 4276 52796
rect 4300 52794 4356 52796
rect 4380 52794 4436 52796
rect 4460 52794 4516 52796
rect 4220 52742 4266 52794
rect 4266 52742 4276 52794
rect 4300 52742 4330 52794
rect 4330 52742 4342 52794
rect 4342 52742 4356 52794
rect 4380 52742 4394 52794
rect 4394 52742 4406 52794
rect 4406 52742 4436 52794
rect 4460 52742 4470 52794
rect 4470 52742 4516 52794
rect 4220 52740 4276 52742
rect 4300 52740 4356 52742
rect 4380 52740 4436 52742
rect 4460 52740 4516 52742
rect 4220 51706 4276 51708
rect 4300 51706 4356 51708
rect 4380 51706 4436 51708
rect 4460 51706 4516 51708
rect 4220 51654 4266 51706
rect 4266 51654 4276 51706
rect 4300 51654 4330 51706
rect 4330 51654 4342 51706
rect 4342 51654 4356 51706
rect 4380 51654 4394 51706
rect 4394 51654 4406 51706
rect 4406 51654 4436 51706
rect 4460 51654 4470 51706
rect 4470 51654 4516 51706
rect 4220 51652 4276 51654
rect 4300 51652 4356 51654
rect 4380 51652 4436 51654
rect 4460 51652 4516 51654
rect 4220 50618 4276 50620
rect 4300 50618 4356 50620
rect 4380 50618 4436 50620
rect 4460 50618 4516 50620
rect 4220 50566 4266 50618
rect 4266 50566 4276 50618
rect 4300 50566 4330 50618
rect 4330 50566 4342 50618
rect 4342 50566 4356 50618
rect 4380 50566 4394 50618
rect 4394 50566 4406 50618
rect 4406 50566 4436 50618
rect 4460 50566 4470 50618
rect 4470 50566 4516 50618
rect 4220 50564 4276 50566
rect 4300 50564 4356 50566
rect 4380 50564 4436 50566
rect 4460 50564 4516 50566
rect 2778 50360 2834 50416
rect 4220 49530 4276 49532
rect 4300 49530 4356 49532
rect 4380 49530 4436 49532
rect 4460 49530 4516 49532
rect 4220 49478 4266 49530
rect 4266 49478 4276 49530
rect 4300 49478 4330 49530
rect 4330 49478 4342 49530
rect 4342 49478 4356 49530
rect 4380 49478 4394 49530
rect 4394 49478 4406 49530
rect 4406 49478 4436 49530
rect 4460 49478 4470 49530
rect 4470 49478 4516 49530
rect 4220 49476 4276 49478
rect 4300 49476 4356 49478
rect 4380 49476 4436 49478
rect 4460 49476 4516 49478
rect 4220 48442 4276 48444
rect 4300 48442 4356 48444
rect 4380 48442 4436 48444
rect 4460 48442 4516 48444
rect 4220 48390 4266 48442
rect 4266 48390 4276 48442
rect 4300 48390 4330 48442
rect 4330 48390 4342 48442
rect 4342 48390 4356 48442
rect 4380 48390 4394 48442
rect 4394 48390 4406 48442
rect 4406 48390 4436 48442
rect 4460 48390 4470 48442
rect 4470 48390 4516 48442
rect 4220 48388 4276 48390
rect 4300 48388 4356 48390
rect 4380 48388 4436 48390
rect 4460 48388 4516 48390
rect 2778 47640 2834 47696
rect 4220 47354 4276 47356
rect 4300 47354 4356 47356
rect 4380 47354 4436 47356
rect 4460 47354 4516 47356
rect 4220 47302 4266 47354
rect 4266 47302 4276 47354
rect 4300 47302 4330 47354
rect 4330 47302 4342 47354
rect 4342 47302 4356 47354
rect 4380 47302 4394 47354
rect 4394 47302 4406 47354
rect 4406 47302 4436 47354
rect 4460 47302 4470 47354
rect 4470 47302 4516 47354
rect 4220 47300 4276 47302
rect 4300 47300 4356 47302
rect 4380 47300 4436 47302
rect 4460 47300 4516 47302
rect 4220 46266 4276 46268
rect 4300 46266 4356 46268
rect 4380 46266 4436 46268
rect 4460 46266 4516 46268
rect 4220 46214 4266 46266
rect 4266 46214 4276 46266
rect 4300 46214 4330 46266
rect 4330 46214 4342 46266
rect 4342 46214 4356 46266
rect 4380 46214 4394 46266
rect 4394 46214 4406 46266
rect 4406 46214 4436 46266
rect 4460 46214 4470 46266
rect 4470 46214 4516 46266
rect 4220 46212 4276 46214
rect 4300 46212 4356 46214
rect 4380 46212 4436 46214
rect 4460 46212 4516 46214
rect 4220 45178 4276 45180
rect 4300 45178 4356 45180
rect 4380 45178 4436 45180
rect 4460 45178 4516 45180
rect 4220 45126 4266 45178
rect 4266 45126 4276 45178
rect 4300 45126 4330 45178
rect 4330 45126 4342 45178
rect 4342 45126 4356 45178
rect 4380 45126 4394 45178
rect 4394 45126 4406 45178
rect 4406 45126 4436 45178
rect 4460 45126 4470 45178
rect 4470 45126 4516 45178
rect 4220 45124 4276 45126
rect 4300 45124 4356 45126
rect 4380 45124 4436 45126
rect 4460 45124 4516 45126
rect 2778 44920 2834 44976
rect 2134 34720 2190 34776
rect 4220 44090 4276 44092
rect 4300 44090 4356 44092
rect 4380 44090 4436 44092
rect 4460 44090 4516 44092
rect 4220 44038 4266 44090
rect 4266 44038 4276 44090
rect 4300 44038 4330 44090
rect 4330 44038 4342 44090
rect 4342 44038 4356 44090
rect 4380 44038 4394 44090
rect 4394 44038 4406 44090
rect 4406 44038 4436 44090
rect 4460 44038 4470 44090
rect 4470 44038 4516 44090
rect 4220 44036 4276 44038
rect 4300 44036 4356 44038
rect 4380 44036 4436 44038
rect 4460 44036 4516 44038
rect 2778 42880 2834 42936
rect 4220 43002 4276 43004
rect 4300 43002 4356 43004
rect 4380 43002 4436 43004
rect 4460 43002 4516 43004
rect 4220 42950 4266 43002
rect 4266 42950 4276 43002
rect 4300 42950 4330 43002
rect 4330 42950 4342 43002
rect 4342 42950 4356 43002
rect 4380 42950 4394 43002
rect 4394 42950 4406 43002
rect 4406 42950 4436 43002
rect 4460 42950 4470 43002
rect 4470 42950 4516 43002
rect 4220 42948 4276 42950
rect 4300 42948 4356 42950
rect 4380 42948 4436 42950
rect 4460 42948 4516 42950
rect 4220 41914 4276 41916
rect 4300 41914 4356 41916
rect 4380 41914 4436 41916
rect 4460 41914 4516 41916
rect 4220 41862 4266 41914
rect 4266 41862 4276 41914
rect 4300 41862 4330 41914
rect 4330 41862 4342 41914
rect 4342 41862 4356 41914
rect 4380 41862 4394 41914
rect 4394 41862 4406 41914
rect 4406 41862 4436 41914
rect 4460 41862 4470 41914
rect 4470 41862 4516 41914
rect 4220 41860 4276 41862
rect 4300 41860 4356 41862
rect 4380 41860 4436 41862
rect 4460 41860 4516 41862
rect 4220 40826 4276 40828
rect 4300 40826 4356 40828
rect 4380 40826 4436 40828
rect 4460 40826 4516 40828
rect 4220 40774 4266 40826
rect 4266 40774 4276 40826
rect 4300 40774 4330 40826
rect 4330 40774 4342 40826
rect 4342 40774 4356 40826
rect 4380 40774 4394 40826
rect 4394 40774 4406 40826
rect 4406 40774 4436 40826
rect 4460 40774 4470 40826
rect 4470 40774 4516 40826
rect 4220 40772 4276 40774
rect 4300 40772 4356 40774
rect 4380 40772 4436 40774
rect 4460 40772 4516 40774
rect 4220 39738 4276 39740
rect 4300 39738 4356 39740
rect 4380 39738 4436 39740
rect 4460 39738 4516 39740
rect 4220 39686 4266 39738
rect 4266 39686 4276 39738
rect 4300 39686 4330 39738
rect 4330 39686 4342 39738
rect 4342 39686 4356 39738
rect 4380 39686 4394 39738
rect 4394 39686 4406 39738
rect 4406 39686 4436 39738
rect 4460 39686 4470 39738
rect 4470 39686 4516 39738
rect 4220 39684 4276 39686
rect 4300 39684 4356 39686
rect 4380 39684 4436 39686
rect 4460 39684 4516 39686
rect 4220 38650 4276 38652
rect 4300 38650 4356 38652
rect 4380 38650 4436 38652
rect 4460 38650 4516 38652
rect 4220 38598 4266 38650
rect 4266 38598 4276 38650
rect 4300 38598 4330 38650
rect 4330 38598 4342 38650
rect 4342 38598 4356 38650
rect 4380 38598 4394 38650
rect 4394 38598 4406 38650
rect 4406 38598 4436 38650
rect 4460 38598 4470 38650
rect 4470 38598 4516 38650
rect 4220 38596 4276 38598
rect 4300 38596 4356 38598
rect 4380 38596 4436 38598
rect 4460 38596 4516 38598
rect 4220 37562 4276 37564
rect 4300 37562 4356 37564
rect 4380 37562 4436 37564
rect 4460 37562 4516 37564
rect 4220 37510 4266 37562
rect 4266 37510 4276 37562
rect 4300 37510 4330 37562
rect 4330 37510 4342 37562
rect 4342 37510 4356 37562
rect 4380 37510 4394 37562
rect 4394 37510 4406 37562
rect 4406 37510 4436 37562
rect 4460 37510 4470 37562
rect 4470 37510 4516 37562
rect 4220 37508 4276 37510
rect 4300 37508 4356 37510
rect 4380 37508 4436 37510
rect 4460 37508 4516 37510
rect 4220 36474 4276 36476
rect 4300 36474 4356 36476
rect 4380 36474 4436 36476
rect 4460 36474 4516 36476
rect 4220 36422 4266 36474
rect 4266 36422 4276 36474
rect 4300 36422 4330 36474
rect 4330 36422 4342 36474
rect 4342 36422 4356 36474
rect 4380 36422 4394 36474
rect 4394 36422 4406 36474
rect 4406 36422 4436 36474
rect 4460 36422 4470 36474
rect 4470 36422 4516 36474
rect 4220 36420 4276 36422
rect 4300 36420 4356 36422
rect 4380 36420 4436 36422
rect 4460 36420 4516 36422
rect 4220 35386 4276 35388
rect 4300 35386 4356 35388
rect 4380 35386 4436 35388
rect 4460 35386 4516 35388
rect 4220 35334 4266 35386
rect 4266 35334 4276 35386
rect 4300 35334 4330 35386
rect 4330 35334 4342 35386
rect 4342 35334 4356 35386
rect 4380 35334 4394 35386
rect 4394 35334 4406 35386
rect 4406 35334 4436 35386
rect 4460 35334 4470 35386
rect 4470 35334 4516 35386
rect 4220 35332 4276 35334
rect 4300 35332 4356 35334
rect 4380 35332 4436 35334
rect 4460 35332 4516 35334
rect 4220 34298 4276 34300
rect 4300 34298 4356 34300
rect 4380 34298 4436 34300
rect 4460 34298 4516 34300
rect 4220 34246 4266 34298
rect 4266 34246 4276 34298
rect 4300 34246 4330 34298
rect 4330 34246 4342 34298
rect 4342 34246 4356 34298
rect 4380 34246 4394 34298
rect 4394 34246 4406 34298
rect 4406 34246 4436 34298
rect 4460 34246 4470 34298
rect 4470 34246 4516 34298
rect 4220 34244 4276 34246
rect 4300 34244 4356 34246
rect 4380 34244 4436 34246
rect 4460 34244 4516 34246
rect 4220 33210 4276 33212
rect 4300 33210 4356 33212
rect 4380 33210 4436 33212
rect 4460 33210 4516 33212
rect 4220 33158 4266 33210
rect 4266 33158 4276 33210
rect 4300 33158 4330 33210
rect 4330 33158 4342 33210
rect 4342 33158 4356 33210
rect 4380 33158 4394 33210
rect 4394 33158 4406 33210
rect 4406 33158 4436 33210
rect 4460 33158 4470 33210
rect 4470 33158 4516 33210
rect 4220 33156 4276 33158
rect 4300 33156 4356 33158
rect 4380 33156 4436 33158
rect 4460 33156 4516 33158
rect 4220 32122 4276 32124
rect 4300 32122 4356 32124
rect 4380 32122 4436 32124
rect 4460 32122 4516 32124
rect 4220 32070 4266 32122
rect 4266 32070 4276 32122
rect 4300 32070 4330 32122
rect 4330 32070 4342 32122
rect 4342 32070 4356 32122
rect 4380 32070 4394 32122
rect 4394 32070 4406 32122
rect 4406 32070 4436 32122
rect 4460 32070 4470 32122
rect 4470 32070 4516 32122
rect 4220 32068 4276 32070
rect 4300 32068 4356 32070
rect 4380 32068 4436 32070
rect 4460 32068 4516 32070
rect 4220 31034 4276 31036
rect 4300 31034 4356 31036
rect 4380 31034 4436 31036
rect 4460 31034 4516 31036
rect 4220 30982 4266 31034
rect 4266 30982 4276 31034
rect 4300 30982 4330 31034
rect 4330 30982 4342 31034
rect 4342 30982 4356 31034
rect 4380 30982 4394 31034
rect 4394 30982 4406 31034
rect 4406 30982 4436 31034
rect 4460 30982 4470 31034
rect 4470 30982 4516 31034
rect 4220 30980 4276 30982
rect 4300 30980 4356 30982
rect 4380 30980 4436 30982
rect 4460 30980 4516 30982
rect 4220 29946 4276 29948
rect 4300 29946 4356 29948
rect 4380 29946 4436 29948
rect 4460 29946 4516 29948
rect 4220 29894 4266 29946
rect 4266 29894 4276 29946
rect 4300 29894 4330 29946
rect 4330 29894 4342 29946
rect 4342 29894 4356 29946
rect 4380 29894 4394 29946
rect 4394 29894 4406 29946
rect 4406 29894 4436 29946
rect 4460 29894 4470 29946
rect 4470 29894 4516 29946
rect 4220 29892 4276 29894
rect 4300 29892 4356 29894
rect 4380 29892 4436 29894
rect 4460 29892 4516 29894
rect 4220 28858 4276 28860
rect 4300 28858 4356 28860
rect 4380 28858 4436 28860
rect 4460 28858 4516 28860
rect 4220 28806 4266 28858
rect 4266 28806 4276 28858
rect 4300 28806 4330 28858
rect 4330 28806 4342 28858
rect 4342 28806 4356 28858
rect 4380 28806 4394 28858
rect 4394 28806 4406 28858
rect 4406 28806 4436 28858
rect 4460 28806 4470 28858
rect 4470 28806 4516 28858
rect 4220 28804 4276 28806
rect 4300 28804 4356 28806
rect 4380 28804 4436 28806
rect 4460 28804 4516 28806
rect 4220 27770 4276 27772
rect 4300 27770 4356 27772
rect 4380 27770 4436 27772
rect 4460 27770 4516 27772
rect 4220 27718 4266 27770
rect 4266 27718 4276 27770
rect 4300 27718 4330 27770
rect 4330 27718 4342 27770
rect 4342 27718 4356 27770
rect 4380 27718 4394 27770
rect 4394 27718 4406 27770
rect 4406 27718 4436 27770
rect 4460 27718 4470 27770
rect 4470 27718 4516 27770
rect 4220 27716 4276 27718
rect 4300 27716 4356 27718
rect 4380 27716 4436 27718
rect 4460 27716 4516 27718
rect 4220 26682 4276 26684
rect 4300 26682 4356 26684
rect 4380 26682 4436 26684
rect 4460 26682 4516 26684
rect 4220 26630 4266 26682
rect 4266 26630 4276 26682
rect 4300 26630 4330 26682
rect 4330 26630 4342 26682
rect 4342 26630 4356 26682
rect 4380 26630 4394 26682
rect 4394 26630 4406 26682
rect 4406 26630 4436 26682
rect 4460 26630 4470 26682
rect 4470 26630 4516 26682
rect 4220 26628 4276 26630
rect 4300 26628 4356 26630
rect 4380 26628 4436 26630
rect 4460 26628 4516 26630
rect 4220 25594 4276 25596
rect 4300 25594 4356 25596
rect 4380 25594 4436 25596
rect 4460 25594 4516 25596
rect 4220 25542 4266 25594
rect 4266 25542 4276 25594
rect 4300 25542 4330 25594
rect 4330 25542 4342 25594
rect 4342 25542 4356 25594
rect 4380 25542 4394 25594
rect 4394 25542 4406 25594
rect 4406 25542 4436 25594
rect 4460 25542 4470 25594
rect 4470 25542 4516 25594
rect 4220 25540 4276 25542
rect 4300 25540 4356 25542
rect 4380 25540 4436 25542
rect 4460 25540 4516 25542
rect 4220 24506 4276 24508
rect 4300 24506 4356 24508
rect 4380 24506 4436 24508
rect 4460 24506 4516 24508
rect 4220 24454 4266 24506
rect 4266 24454 4276 24506
rect 4300 24454 4330 24506
rect 4330 24454 4342 24506
rect 4342 24454 4356 24506
rect 4380 24454 4394 24506
rect 4394 24454 4406 24506
rect 4406 24454 4436 24506
rect 4460 24454 4470 24506
rect 4470 24454 4516 24506
rect 4220 24452 4276 24454
rect 4300 24452 4356 24454
rect 4380 24452 4436 24454
rect 4460 24452 4516 24454
rect 4220 23418 4276 23420
rect 4300 23418 4356 23420
rect 4380 23418 4436 23420
rect 4460 23418 4516 23420
rect 4220 23366 4266 23418
rect 4266 23366 4276 23418
rect 4300 23366 4330 23418
rect 4330 23366 4342 23418
rect 4342 23366 4356 23418
rect 4380 23366 4394 23418
rect 4394 23366 4406 23418
rect 4406 23366 4436 23418
rect 4460 23366 4470 23418
rect 4470 23366 4516 23418
rect 4220 23364 4276 23366
rect 4300 23364 4356 23366
rect 4380 23364 4436 23366
rect 4460 23364 4516 23366
rect 4220 22330 4276 22332
rect 4300 22330 4356 22332
rect 4380 22330 4436 22332
rect 4460 22330 4516 22332
rect 4220 22278 4266 22330
rect 4266 22278 4276 22330
rect 4300 22278 4330 22330
rect 4330 22278 4342 22330
rect 4342 22278 4356 22330
rect 4380 22278 4394 22330
rect 4394 22278 4406 22330
rect 4406 22278 4436 22330
rect 4460 22278 4470 22330
rect 4470 22278 4516 22330
rect 4220 22276 4276 22278
rect 4300 22276 4356 22278
rect 4380 22276 4436 22278
rect 4460 22276 4516 22278
rect 4220 21242 4276 21244
rect 4300 21242 4356 21244
rect 4380 21242 4436 21244
rect 4460 21242 4516 21244
rect 4220 21190 4266 21242
rect 4266 21190 4276 21242
rect 4300 21190 4330 21242
rect 4330 21190 4342 21242
rect 4342 21190 4356 21242
rect 4380 21190 4394 21242
rect 4394 21190 4406 21242
rect 4406 21190 4436 21242
rect 4460 21190 4470 21242
rect 4470 21190 4516 21242
rect 4220 21188 4276 21190
rect 4300 21188 4356 21190
rect 4380 21188 4436 21190
rect 4460 21188 4516 21190
rect 4220 20154 4276 20156
rect 4300 20154 4356 20156
rect 4380 20154 4436 20156
rect 4460 20154 4516 20156
rect 4220 20102 4266 20154
rect 4266 20102 4276 20154
rect 4300 20102 4330 20154
rect 4330 20102 4342 20154
rect 4342 20102 4356 20154
rect 4380 20102 4394 20154
rect 4394 20102 4406 20154
rect 4406 20102 4436 20154
rect 4460 20102 4470 20154
rect 4470 20102 4516 20154
rect 4220 20100 4276 20102
rect 4300 20100 4356 20102
rect 4380 20100 4436 20102
rect 4460 20100 4516 20102
rect 4220 19066 4276 19068
rect 4300 19066 4356 19068
rect 4380 19066 4436 19068
rect 4460 19066 4516 19068
rect 4220 19014 4266 19066
rect 4266 19014 4276 19066
rect 4300 19014 4330 19066
rect 4330 19014 4342 19066
rect 4342 19014 4356 19066
rect 4380 19014 4394 19066
rect 4394 19014 4406 19066
rect 4406 19014 4436 19066
rect 4460 19014 4470 19066
rect 4470 19014 4516 19066
rect 4220 19012 4276 19014
rect 4300 19012 4356 19014
rect 4380 19012 4436 19014
rect 4460 19012 4516 19014
rect 4220 17978 4276 17980
rect 4300 17978 4356 17980
rect 4380 17978 4436 17980
rect 4460 17978 4516 17980
rect 4220 17926 4266 17978
rect 4266 17926 4276 17978
rect 4300 17926 4330 17978
rect 4330 17926 4342 17978
rect 4342 17926 4356 17978
rect 4380 17926 4394 17978
rect 4394 17926 4406 17978
rect 4406 17926 4436 17978
rect 4460 17926 4470 17978
rect 4470 17926 4516 17978
rect 4220 17924 4276 17926
rect 4300 17924 4356 17926
rect 4380 17924 4436 17926
rect 4460 17924 4516 17926
rect 4220 16890 4276 16892
rect 4300 16890 4356 16892
rect 4380 16890 4436 16892
rect 4460 16890 4516 16892
rect 4220 16838 4266 16890
rect 4266 16838 4276 16890
rect 4300 16838 4330 16890
rect 4330 16838 4342 16890
rect 4342 16838 4356 16890
rect 4380 16838 4394 16890
rect 4394 16838 4406 16890
rect 4406 16838 4436 16890
rect 4460 16838 4470 16890
rect 4470 16838 4516 16890
rect 4220 16836 4276 16838
rect 4300 16836 4356 16838
rect 4380 16836 4436 16838
rect 4460 16836 4516 16838
rect 19580 55514 19636 55516
rect 19660 55514 19716 55516
rect 19740 55514 19796 55516
rect 19820 55514 19876 55516
rect 19580 55462 19626 55514
rect 19626 55462 19636 55514
rect 19660 55462 19690 55514
rect 19690 55462 19702 55514
rect 19702 55462 19716 55514
rect 19740 55462 19754 55514
rect 19754 55462 19766 55514
rect 19766 55462 19796 55514
rect 19820 55462 19830 55514
rect 19830 55462 19876 55514
rect 19580 55460 19636 55462
rect 19660 55460 19716 55462
rect 19740 55460 19796 55462
rect 19820 55460 19876 55462
rect 34940 57146 34996 57148
rect 35020 57146 35076 57148
rect 35100 57146 35156 57148
rect 35180 57146 35236 57148
rect 34940 57094 34986 57146
rect 34986 57094 34996 57146
rect 35020 57094 35050 57146
rect 35050 57094 35062 57146
rect 35062 57094 35076 57146
rect 35100 57094 35114 57146
rect 35114 57094 35126 57146
rect 35126 57094 35156 57146
rect 35180 57094 35190 57146
rect 35190 57094 35236 57146
rect 34940 57092 34996 57094
rect 35020 57092 35076 57094
rect 35100 57092 35156 57094
rect 35180 57092 35236 57094
rect 34940 56058 34996 56060
rect 35020 56058 35076 56060
rect 35100 56058 35156 56060
rect 35180 56058 35236 56060
rect 34940 56006 34986 56058
rect 34986 56006 34996 56058
rect 35020 56006 35050 56058
rect 35050 56006 35062 56058
rect 35062 56006 35076 56058
rect 35100 56006 35114 56058
rect 35114 56006 35126 56058
rect 35126 56006 35156 56058
rect 35180 56006 35190 56058
rect 35190 56006 35236 56058
rect 34940 56004 34996 56006
rect 35020 56004 35076 56006
rect 35100 56004 35156 56006
rect 35180 56004 35236 56006
rect 50300 57690 50356 57692
rect 50380 57690 50436 57692
rect 50460 57690 50516 57692
rect 50540 57690 50596 57692
rect 50300 57638 50346 57690
rect 50346 57638 50356 57690
rect 50380 57638 50410 57690
rect 50410 57638 50422 57690
rect 50422 57638 50436 57690
rect 50460 57638 50474 57690
rect 50474 57638 50486 57690
rect 50486 57638 50516 57690
rect 50540 57638 50550 57690
rect 50550 57638 50596 57690
rect 50300 57636 50356 57638
rect 50380 57636 50436 57638
rect 50460 57636 50516 57638
rect 50540 57636 50596 57638
rect 4220 15802 4276 15804
rect 4300 15802 4356 15804
rect 4380 15802 4436 15804
rect 4460 15802 4516 15804
rect 4220 15750 4266 15802
rect 4266 15750 4276 15802
rect 4300 15750 4330 15802
rect 4330 15750 4342 15802
rect 4342 15750 4356 15802
rect 4380 15750 4394 15802
rect 4394 15750 4406 15802
rect 4406 15750 4436 15802
rect 4460 15750 4470 15802
rect 4470 15750 4516 15802
rect 4220 15748 4276 15750
rect 4300 15748 4356 15750
rect 4380 15748 4436 15750
rect 4460 15748 4516 15750
rect 4220 14714 4276 14716
rect 4300 14714 4356 14716
rect 4380 14714 4436 14716
rect 4460 14714 4516 14716
rect 4220 14662 4266 14714
rect 4266 14662 4276 14714
rect 4300 14662 4330 14714
rect 4330 14662 4342 14714
rect 4342 14662 4356 14714
rect 4380 14662 4394 14714
rect 4394 14662 4406 14714
rect 4406 14662 4436 14714
rect 4460 14662 4470 14714
rect 4470 14662 4516 14714
rect 4220 14660 4276 14662
rect 4300 14660 4356 14662
rect 4380 14660 4436 14662
rect 4460 14660 4516 14662
rect 4220 13626 4276 13628
rect 4300 13626 4356 13628
rect 4380 13626 4436 13628
rect 4460 13626 4516 13628
rect 4220 13574 4266 13626
rect 4266 13574 4276 13626
rect 4300 13574 4330 13626
rect 4330 13574 4342 13626
rect 4342 13574 4356 13626
rect 4380 13574 4394 13626
rect 4394 13574 4406 13626
rect 4406 13574 4436 13626
rect 4460 13574 4470 13626
rect 4470 13574 4516 13626
rect 4220 13572 4276 13574
rect 4300 13572 4356 13574
rect 4380 13572 4436 13574
rect 4460 13572 4516 13574
rect 4220 12538 4276 12540
rect 4300 12538 4356 12540
rect 4380 12538 4436 12540
rect 4460 12538 4516 12540
rect 4220 12486 4266 12538
rect 4266 12486 4276 12538
rect 4300 12486 4330 12538
rect 4330 12486 4342 12538
rect 4342 12486 4356 12538
rect 4380 12486 4394 12538
rect 4394 12486 4406 12538
rect 4406 12486 4436 12538
rect 4460 12486 4470 12538
rect 4470 12486 4516 12538
rect 4220 12484 4276 12486
rect 4300 12484 4356 12486
rect 4380 12484 4436 12486
rect 4460 12484 4516 12486
rect 4220 11450 4276 11452
rect 4300 11450 4356 11452
rect 4380 11450 4436 11452
rect 4460 11450 4516 11452
rect 4220 11398 4266 11450
rect 4266 11398 4276 11450
rect 4300 11398 4330 11450
rect 4330 11398 4342 11450
rect 4342 11398 4356 11450
rect 4380 11398 4394 11450
rect 4394 11398 4406 11450
rect 4406 11398 4436 11450
rect 4460 11398 4470 11450
rect 4470 11398 4516 11450
rect 4220 11396 4276 11398
rect 4300 11396 4356 11398
rect 4380 11396 4436 11398
rect 4460 11396 4516 11398
rect 4220 10362 4276 10364
rect 4300 10362 4356 10364
rect 4380 10362 4436 10364
rect 4460 10362 4516 10364
rect 4220 10310 4266 10362
rect 4266 10310 4276 10362
rect 4300 10310 4330 10362
rect 4330 10310 4342 10362
rect 4342 10310 4356 10362
rect 4380 10310 4394 10362
rect 4394 10310 4406 10362
rect 4406 10310 4436 10362
rect 4460 10310 4470 10362
rect 4470 10310 4516 10362
rect 4220 10308 4276 10310
rect 4300 10308 4356 10310
rect 4380 10308 4436 10310
rect 4460 10308 4516 10310
rect 2778 9560 2834 9616
rect 4220 9274 4276 9276
rect 4300 9274 4356 9276
rect 4380 9274 4436 9276
rect 4460 9274 4516 9276
rect 4220 9222 4266 9274
rect 4266 9222 4276 9274
rect 4300 9222 4330 9274
rect 4330 9222 4342 9274
rect 4342 9222 4356 9274
rect 4380 9222 4394 9274
rect 4394 9222 4406 9274
rect 4406 9222 4436 9274
rect 4460 9222 4470 9274
rect 4470 9222 4516 9274
rect 4220 9220 4276 9222
rect 4300 9220 4356 9222
rect 4380 9220 4436 9222
rect 4460 9220 4516 9222
rect 4220 8186 4276 8188
rect 4300 8186 4356 8188
rect 4380 8186 4436 8188
rect 4460 8186 4516 8188
rect 4220 8134 4266 8186
rect 4266 8134 4276 8186
rect 4300 8134 4330 8186
rect 4330 8134 4342 8186
rect 4342 8134 4356 8186
rect 4380 8134 4394 8186
rect 4394 8134 4406 8186
rect 4406 8134 4436 8186
rect 4460 8134 4470 8186
rect 4470 8134 4516 8186
rect 4220 8132 4276 8134
rect 4300 8132 4356 8134
rect 4380 8132 4436 8134
rect 4460 8132 4516 8134
rect 4220 7098 4276 7100
rect 4300 7098 4356 7100
rect 4380 7098 4436 7100
rect 4460 7098 4516 7100
rect 4220 7046 4266 7098
rect 4266 7046 4276 7098
rect 4300 7046 4330 7098
rect 4330 7046 4342 7098
rect 4342 7046 4356 7098
rect 4380 7046 4394 7098
rect 4394 7046 4406 7098
rect 4406 7046 4436 7098
rect 4460 7046 4470 7098
rect 4470 7046 4516 7098
rect 4220 7044 4276 7046
rect 4300 7044 4356 7046
rect 4380 7044 4436 7046
rect 4460 7044 4516 7046
rect 4220 6010 4276 6012
rect 4300 6010 4356 6012
rect 4380 6010 4436 6012
rect 4460 6010 4516 6012
rect 4220 5958 4266 6010
rect 4266 5958 4276 6010
rect 4300 5958 4330 6010
rect 4330 5958 4342 6010
rect 4342 5958 4356 6010
rect 4380 5958 4394 6010
rect 4394 5958 4406 6010
rect 4406 5958 4436 6010
rect 4460 5958 4470 6010
rect 4470 5958 4516 6010
rect 4220 5956 4276 5958
rect 4300 5956 4356 5958
rect 4380 5956 4436 5958
rect 4460 5956 4516 5958
rect 4220 4922 4276 4924
rect 4300 4922 4356 4924
rect 4380 4922 4436 4924
rect 4460 4922 4516 4924
rect 4220 4870 4266 4922
rect 4266 4870 4276 4922
rect 4300 4870 4330 4922
rect 4330 4870 4342 4922
rect 4342 4870 4356 4922
rect 4380 4870 4394 4922
rect 4394 4870 4406 4922
rect 4406 4870 4436 4922
rect 4460 4870 4470 4922
rect 4470 4870 4516 4922
rect 4220 4868 4276 4870
rect 4300 4868 4356 4870
rect 4380 4868 4436 4870
rect 4460 4868 4516 4870
rect 2778 4800 2834 4856
rect 19580 54426 19636 54428
rect 19660 54426 19716 54428
rect 19740 54426 19796 54428
rect 19820 54426 19876 54428
rect 19580 54374 19626 54426
rect 19626 54374 19636 54426
rect 19660 54374 19690 54426
rect 19690 54374 19702 54426
rect 19702 54374 19716 54426
rect 19740 54374 19754 54426
rect 19754 54374 19766 54426
rect 19766 54374 19796 54426
rect 19820 54374 19830 54426
rect 19830 54374 19876 54426
rect 19580 54372 19636 54374
rect 19660 54372 19716 54374
rect 19740 54372 19796 54374
rect 19820 54372 19876 54374
rect 19580 53338 19636 53340
rect 19660 53338 19716 53340
rect 19740 53338 19796 53340
rect 19820 53338 19876 53340
rect 19580 53286 19626 53338
rect 19626 53286 19636 53338
rect 19660 53286 19690 53338
rect 19690 53286 19702 53338
rect 19702 53286 19716 53338
rect 19740 53286 19754 53338
rect 19754 53286 19766 53338
rect 19766 53286 19796 53338
rect 19820 53286 19830 53338
rect 19830 53286 19876 53338
rect 19580 53284 19636 53286
rect 19660 53284 19716 53286
rect 19740 53284 19796 53286
rect 19820 53284 19876 53286
rect 19580 52250 19636 52252
rect 19660 52250 19716 52252
rect 19740 52250 19796 52252
rect 19820 52250 19876 52252
rect 19580 52198 19626 52250
rect 19626 52198 19636 52250
rect 19660 52198 19690 52250
rect 19690 52198 19702 52250
rect 19702 52198 19716 52250
rect 19740 52198 19754 52250
rect 19754 52198 19766 52250
rect 19766 52198 19796 52250
rect 19820 52198 19830 52250
rect 19830 52198 19876 52250
rect 19580 52196 19636 52198
rect 19660 52196 19716 52198
rect 19740 52196 19796 52198
rect 19820 52196 19876 52198
rect 19580 51162 19636 51164
rect 19660 51162 19716 51164
rect 19740 51162 19796 51164
rect 19820 51162 19876 51164
rect 19580 51110 19626 51162
rect 19626 51110 19636 51162
rect 19660 51110 19690 51162
rect 19690 51110 19702 51162
rect 19702 51110 19716 51162
rect 19740 51110 19754 51162
rect 19754 51110 19766 51162
rect 19766 51110 19796 51162
rect 19820 51110 19830 51162
rect 19830 51110 19876 51162
rect 19580 51108 19636 51110
rect 19660 51108 19716 51110
rect 19740 51108 19796 51110
rect 19820 51108 19876 51110
rect 19580 50074 19636 50076
rect 19660 50074 19716 50076
rect 19740 50074 19796 50076
rect 19820 50074 19876 50076
rect 19580 50022 19626 50074
rect 19626 50022 19636 50074
rect 19660 50022 19690 50074
rect 19690 50022 19702 50074
rect 19702 50022 19716 50074
rect 19740 50022 19754 50074
rect 19754 50022 19766 50074
rect 19766 50022 19796 50074
rect 19820 50022 19830 50074
rect 19830 50022 19876 50074
rect 19580 50020 19636 50022
rect 19660 50020 19716 50022
rect 19740 50020 19796 50022
rect 19820 50020 19876 50022
rect 19580 48986 19636 48988
rect 19660 48986 19716 48988
rect 19740 48986 19796 48988
rect 19820 48986 19876 48988
rect 19580 48934 19626 48986
rect 19626 48934 19636 48986
rect 19660 48934 19690 48986
rect 19690 48934 19702 48986
rect 19702 48934 19716 48986
rect 19740 48934 19754 48986
rect 19754 48934 19766 48986
rect 19766 48934 19796 48986
rect 19820 48934 19830 48986
rect 19830 48934 19876 48986
rect 19580 48932 19636 48934
rect 19660 48932 19716 48934
rect 19740 48932 19796 48934
rect 19820 48932 19876 48934
rect 19580 47898 19636 47900
rect 19660 47898 19716 47900
rect 19740 47898 19796 47900
rect 19820 47898 19876 47900
rect 19580 47846 19626 47898
rect 19626 47846 19636 47898
rect 19660 47846 19690 47898
rect 19690 47846 19702 47898
rect 19702 47846 19716 47898
rect 19740 47846 19754 47898
rect 19754 47846 19766 47898
rect 19766 47846 19796 47898
rect 19820 47846 19830 47898
rect 19830 47846 19876 47898
rect 19580 47844 19636 47846
rect 19660 47844 19716 47846
rect 19740 47844 19796 47846
rect 19820 47844 19876 47846
rect 19580 46810 19636 46812
rect 19660 46810 19716 46812
rect 19740 46810 19796 46812
rect 19820 46810 19876 46812
rect 19580 46758 19626 46810
rect 19626 46758 19636 46810
rect 19660 46758 19690 46810
rect 19690 46758 19702 46810
rect 19702 46758 19716 46810
rect 19740 46758 19754 46810
rect 19754 46758 19766 46810
rect 19766 46758 19796 46810
rect 19820 46758 19830 46810
rect 19830 46758 19876 46810
rect 19580 46756 19636 46758
rect 19660 46756 19716 46758
rect 19740 46756 19796 46758
rect 19820 46756 19876 46758
rect 19580 45722 19636 45724
rect 19660 45722 19716 45724
rect 19740 45722 19796 45724
rect 19820 45722 19876 45724
rect 19580 45670 19626 45722
rect 19626 45670 19636 45722
rect 19660 45670 19690 45722
rect 19690 45670 19702 45722
rect 19702 45670 19716 45722
rect 19740 45670 19754 45722
rect 19754 45670 19766 45722
rect 19766 45670 19796 45722
rect 19820 45670 19830 45722
rect 19830 45670 19876 45722
rect 19580 45668 19636 45670
rect 19660 45668 19716 45670
rect 19740 45668 19796 45670
rect 19820 45668 19876 45670
rect 19580 44634 19636 44636
rect 19660 44634 19716 44636
rect 19740 44634 19796 44636
rect 19820 44634 19876 44636
rect 19580 44582 19626 44634
rect 19626 44582 19636 44634
rect 19660 44582 19690 44634
rect 19690 44582 19702 44634
rect 19702 44582 19716 44634
rect 19740 44582 19754 44634
rect 19754 44582 19766 44634
rect 19766 44582 19796 44634
rect 19820 44582 19830 44634
rect 19830 44582 19876 44634
rect 19580 44580 19636 44582
rect 19660 44580 19716 44582
rect 19740 44580 19796 44582
rect 19820 44580 19876 44582
rect 19580 43546 19636 43548
rect 19660 43546 19716 43548
rect 19740 43546 19796 43548
rect 19820 43546 19876 43548
rect 19580 43494 19626 43546
rect 19626 43494 19636 43546
rect 19660 43494 19690 43546
rect 19690 43494 19702 43546
rect 19702 43494 19716 43546
rect 19740 43494 19754 43546
rect 19754 43494 19766 43546
rect 19766 43494 19796 43546
rect 19820 43494 19830 43546
rect 19830 43494 19876 43546
rect 19580 43492 19636 43494
rect 19660 43492 19716 43494
rect 19740 43492 19796 43494
rect 19820 43492 19876 43494
rect 19580 42458 19636 42460
rect 19660 42458 19716 42460
rect 19740 42458 19796 42460
rect 19820 42458 19876 42460
rect 19580 42406 19626 42458
rect 19626 42406 19636 42458
rect 19660 42406 19690 42458
rect 19690 42406 19702 42458
rect 19702 42406 19716 42458
rect 19740 42406 19754 42458
rect 19754 42406 19766 42458
rect 19766 42406 19796 42458
rect 19820 42406 19830 42458
rect 19830 42406 19876 42458
rect 19580 42404 19636 42406
rect 19660 42404 19716 42406
rect 19740 42404 19796 42406
rect 19820 42404 19876 42406
rect 34940 54970 34996 54972
rect 35020 54970 35076 54972
rect 35100 54970 35156 54972
rect 35180 54970 35236 54972
rect 34940 54918 34986 54970
rect 34986 54918 34996 54970
rect 35020 54918 35050 54970
rect 35050 54918 35062 54970
rect 35062 54918 35076 54970
rect 35100 54918 35114 54970
rect 35114 54918 35126 54970
rect 35126 54918 35156 54970
rect 35180 54918 35190 54970
rect 35190 54918 35236 54970
rect 34940 54916 34996 54918
rect 35020 54916 35076 54918
rect 35100 54916 35156 54918
rect 35180 54916 35236 54918
rect 34940 53882 34996 53884
rect 35020 53882 35076 53884
rect 35100 53882 35156 53884
rect 35180 53882 35236 53884
rect 34940 53830 34986 53882
rect 34986 53830 34996 53882
rect 35020 53830 35050 53882
rect 35050 53830 35062 53882
rect 35062 53830 35076 53882
rect 35100 53830 35114 53882
rect 35114 53830 35126 53882
rect 35126 53830 35156 53882
rect 35180 53830 35190 53882
rect 35190 53830 35236 53882
rect 34940 53828 34996 53830
rect 35020 53828 35076 53830
rect 35100 53828 35156 53830
rect 35180 53828 35236 53830
rect 50300 56602 50356 56604
rect 50380 56602 50436 56604
rect 50460 56602 50516 56604
rect 50540 56602 50596 56604
rect 50300 56550 50346 56602
rect 50346 56550 50356 56602
rect 50380 56550 50410 56602
rect 50410 56550 50422 56602
rect 50422 56550 50436 56602
rect 50460 56550 50474 56602
rect 50474 56550 50486 56602
rect 50486 56550 50516 56602
rect 50540 56550 50550 56602
rect 50550 56550 50596 56602
rect 50300 56548 50356 56550
rect 50380 56548 50436 56550
rect 50460 56548 50516 56550
rect 50540 56548 50596 56550
rect 34940 52794 34996 52796
rect 35020 52794 35076 52796
rect 35100 52794 35156 52796
rect 35180 52794 35236 52796
rect 34940 52742 34986 52794
rect 34986 52742 34996 52794
rect 35020 52742 35050 52794
rect 35050 52742 35062 52794
rect 35062 52742 35076 52794
rect 35100 52742 35114 52794
rect 35114 52742 35126 52794
rect 35126 52742 35156 52794
rect 35180 52742 35190 52794
rect 35190 52742 35236 52794
rect 34940 52740 34996 52742
rect 35020 52740 35076 52742
rect 35100 52740 35156 52742
rect 35180 52740 35236 52742
rect 50300 55514 50356 55516
rect 50380 55514 50436 55516
rect 50460 55514 50516 55516
rect 50540 55514 50596 55516
rect 50300 55462 50346 55514
rect 50346 55462 50356 55514
rect 50380 55462 50410 55514
rect 50410 55462 50422 55514
rect 50422 55462 50436 55514
rect 50460 55462 50474 55514
rect 50474 55462 50486 55514
rect 50486 55462 50516 55514
rect 50540 55462 50550 55514
rect 50550 55462 50596 55514
rect 50300 55460 50356 55462
rect 50380 55460 50436 55462
rect 50460 55460 50516 55462
rect 50540 55460 50596 55462
rect 50300 54426 50356 54428
rect 50380 54426 50436 54428
rect 50460 54426 50516 54428
rect 50540 54426 50596 54428
rect 50300 54374 50346 54426
rect 50346 54374 50356 54426
rect 50380 54374 50410 54426
rect 50410 54374 50422 54426
rect 50422 54374 50436 54426
rect 50460 54374 50474 54426
rect 50474 54374 50486 54426
rect 50486 54374 50516 54426
rect 50540 54374 50550 54426
rect 50550 54374 50596 54426
rect 50300 54372 50356 54374
rect 50380 54372 50436 54374
rect 50460 54372 50516 54374
rect 50540 54372 50596 54374
rect 34940 51706 34996 51708
rect 35020 51706 35076 51708
rect 35100 51706 35156 51708
rect 35180 51706 35236 51708
rect 34940 51654 34986 51706
rect 34986 51654 34996 51706
rect 35020 51654 35050 51706
rect 35050 51654 35062 51706
rect 35062 51654 35076 51706
rect 35100 51654 35114 51706
rect 35114 51654 35126 51706
rect 35126 51654 35156 51706
rect 35180 51654 35190 51706
rect 35190 51654 35236 51706
rect 34940 51652 34996 51654
rect 35020 51652 35076 51654
rect 35100 51652 35156 51654
rect 35180 51652 35236 51654
rect 34940 50618 34996 50620
rect 35020 50618 35076 50620
rect 35100 50618 35156 50620
rect 35180 50618 35236 50620
rect 34940 50566 34986 50618
rect 34986 50566 34996 50618
rect 35020 50566 35050 50618
rect 35050 50566 35062 50618
rect 35062 50566 35076 50618
rect 35100 50566 35114 50618
rect 35114 50566 35126 50618
rect 35126 50566 35156 50618
rect 35180 50566 35190 50618
rect 35190 50566 35236 50618
rect 34940 50564 34996 50566
rect 35020 50564 35076 50566
rect 35100 50564 35156 50566
rect 35180 50564 35236 50566
rect 34940 49530 34996 49532
rect 35020 49530 35076 49532
rect 35100 49530 35156 49532
rect 35180 49530 35236 49532
rect 34940 49478 34986 49530
rect 34986 49478 34996 49530
rect 35020 49478 35050 49530
rect 35050 49478 35062 49530
rect 35062 49478 35076 49530
rect 35100 49478 35114 49530
rect 35114 49478 35126 49530
rect 35126 49478 35156 49530
rect 35180 49478 35190 49530
rect 35190 49478 35236 49530
rect 34940 49476 34996 49478
rect 35020 49476 35076 49478
rect 35100 49476 35156 49478
rect 35180 49476 35236 49478
rect 34940 48442 34996 48444
rect 35020 48442 35076 48444
rect 35100 48442 35156 48444
rect 35180 48442 35236 48444
rect 34940 48390 34986 48442
rect 34986 48390 34996 48442
rect 35020 48390 35050 48442
rect 35050 48390 35062 48442
rect 35062 48390 35076 48442
rect 35100 48390 35114 48442
rect 35114 48390 35126 48442
rect 35126 48390 35156 48442
rect 35180 48390 35190 48442
rect 35190 48390 35236 48442
rect 34940 48388 34996 48390
rect 35020 48388 35076 48390
rect 35100 48388 35156 48390
rect 35180 48388 35236 48390
rect 34940 47354 34996 47356
rect 35020 47354 35076 47356
rect 35100 47354 35156 47356
rect 35180 47354 35236 47356
rect 34940 47302 34986 47354
rect 34986 47302 34996 47354
rect 35020 47302 35050 47354
rect 35050 47302 35062 47354
rect 35062 47302 35076 47354
rect 35100 47302 35114 47354
rect 35114 47302 35126 47354
rect 35126 47302 35156 47354
rect 35180 47302 35190 47354
rect 35190 47302 35236 47354
rect 34940 47300 34996 47302
rect 35020 47300 35076 47302
rect 35100 47300 35156 47302
rect 35180 47300 35236 47302
rect 34940 46266 34996 46268
rect 35020 46266 35076 46268
rect 35100 46266 35156 46268
rect 35180 46266 35236 46268
rect 34940 46214 34986 46266
rect 34986 46214 34996 46266
rect 35020 46214 35050 46266
rect 35050 46214 35062 46266
rect 35062 46214 35076 46266
rect 35100 46214 35114 46266
rect 35114 46214 35126 46266
rect 35126 46214 35156 46266
rect 35180 46214 35190 46266
rect 35190 46214 35236 46266
rect 34940 46212 34996 46214
rect 35020 46212 35076 46214
rect 35100 46212 35156 46214
rect 35180 46212 35236 46214
rect 34940 45178 34996 45180
rect 35020 45178 35076 45180
rect 35100 45178 35156 45180
rect 35180 45178 35236 45180
rect 34940 45126 34986 45178
rect 34986 45126 34996 45178
rect 35020 45126 35050 45178
rect 35050 45126 35062 45178
rect 35062 45126 35076 45178
rect 35100 45126 35114 45178
rect 35114 45126 35126 45178
rect 35126 45126 35156 45178
rect 35180 45126 35190 45178
rect 35190 45126 35236 45178
rect 34940 45124 34996 45126
rect 35020 45124 35076 45126
rect 35100 45124 35156 45126
rect 35180 45124 35236 45126
rect 34940 44090 34996 44092
rect 35020 44090 35076 44092
rect 35100 44090 35156 44092
rect 35180 44090 35236 44092
rect 34940 44038 34986 44090
rect 34986 44038 34996 44090
rect 35020 44038 35050 44090
rect 35050 44038 35062 44090
rect 35062 44038 35076 44090
rect 35100 44038 35114 44090
rect 35114 44038 35126 44090
rect 35126 44038 35156 44090
rect 35180 44038 35190 44090
rect 35190 44038 35236 44090
rect 34940 44036 34996 44038
rect 35020 44036 35076 44038
rect 35100 44036 35156 44038
rect 35180 44036 35236 44038
rect 34940 43002 34996 43004
rect 35020 43002 35076 43004
rect 35100 43002 35156 43004
rect 35180 43002 35236 43004
rect 34940 42950 34986 43002
rect 34986 42950 34996 43002
rect 35020 42950 35050 43002
rect 35050 42950 35062 43002
rect 35062 42950 35076 43002
rect 35100 42950 35114 43002
rect 35114 42950 35126 43002
rect 35126 42950 35156 43002
rect 35180 42950 35190 43002
rect 35190 42950 35236 43002
rect 34940 42948 34996 42950
rect 35020 42948 35076 42950
rect 35100 42948 35156 42950
rect 35180 42948 35236 42950
rect 50300 53338 50356 53340
rect 50380 53338 50436 53340
rect 50460 53338 50516 53340
rect 50540 53338 50596 53340
rect 50300 53286 50346 53338
rect 50346 53286 50356 53338
rect 50380 53286 50410 53338
rect 50410 53286 50422 53338
rect 50422 53286 50436 53338
rect 50460 53286 50474 53338
rect 50474 53286 50486 53338
rect 50486 53286 50516 53338
rect 50540 53286 50550 53338
rect 50550 53286 50596 53338
rect 50300 53284 50356 53286
rect 50380 53284 50436 53286
rect 50460 53284 50516 53286
rect 50540 53284 50596 53286
rect 50300 52250 50356 52252
rect 50380 52250 50436 52252
rect 50460 52250 50516 52252
rect 50540 52250 50596 52252
rect 50300 52198 50346 52250
rect 50346 52198 50356 52250
rect 50380 52198 50410 52250
rect 50410 52198 50422 52250
rect 50422 52198 50436 52250
rect 50460 52198 50474 52250
rect 50474 52198 50486 52250
rect 50486 52198 50516 52250
rect 50540 52198 50550 52250
rect 50550 52198 50596 52250
rect 50300 52196 50356 52198
rect 50380 52196 50436 52198
rect 50460 52196 50516 52198
rect 50540 52196 50596 52198
rect 50300 51162 50356 51164
rect 50380 51162 50436 51164
rect 50460 51162 50516 51164
rect 50540 51162 50596 51164
rect 50300 51110 50346 51162
rect 50346 51110 50356 51162
rect 50380 51110 50410 51162
rect 50410 51110 50422 51162
rect 50422 51110 50436 51162
rect 50460 51110 50474 51162
rect 50474 51110 50486 51162
rect 50486 51110 50516 51162
rect 50540 51110 50550 51162
rect 50550 51110 50596 51162
rect 50300 51108 50356 51110
rect 50380 51108 50436 51110
rect 50460 51108 50516 51110
rect 50540 51108 50596 51110
rect 50300 50074 50356 50076
rect 50380 50074 50436 50076
rect 50460 50074 50516 50076
rect 50540 50074 50596 50076
rect 50300 50022 50346 50074
rect 50346 50022 50356 50074
rect 50380 50022 50410 50074
rect 50410 50022 50422 50074
rect 50422 50022 50436 50074
rect 50460 50022 50474 50074
rect 50474 50022 50486 50074
rect 50486 50022 50516 50074
rect 50540 50022 50550 50074
rect 50550 50022 50596 50074
rect 50300 50020 50356 50022
rect 50380 50020 50436 50022
rect 50460 50020 50516 50022
rect 50540 50020 50596 50022
rect 34940 41914 34996 41916
rect 35020 41914 35076 41916
rect 35100 41914 35156 41916
rect 35180 41914 35236 41916
rect 34940 41862 34986 41914
rect 34986 41862 34996 41914
rect 35020 41862 35050 41914
rect 35050 41862 35062 41914
rect 35062 41862 35076 41914
rect 35100 41862 35114 41914
rect 35114 41862 35126 41914
rect 35126 41862 35156 41914
rect 35180 41862 35190 41914
rect 35190 41862 35236 41914
rect 34940 41860 34996 41862
rect 35020 41860 35076 41862
rect 35100 41860 35156 41862
rect 35180 41860 35236 41862
rect 19580 41370 19636 41372
rect 19660 41370 19716 41372
rect 19740 41370 19796 41372
rect 19820 41370 19876 41372
rect 19580 41318 19626 41370
rect 19626 41318 19636 41370
rect 19660 41318 19690 41370
rect 19690 41318 19702 41370
rect 19702 41318 19716 41370
rect 19740 41318 19754 41370
rect 19754 41318 19766 41370
rect 19766 41318 19796 41370
rect 19820 41318 19830 41370
rect 19830 41318 19876 41370
rect 19580 41316 19636 41318
rect 19660 41316 19716 41318
rect 19740 41316 19796 41318
rect 19820 41316 19876 41318
rect 34940 40826 34996 40828
rect 35020 40826 35076 40828
rect 35100 40826 35156 40828
rect 35180 40826 35236 40828
rect 34940 40774 34986 40826
rect 34986 40774 34996 40826
rect 35020 40774 35050 40826
rect 35050 40774 35062 40826
rect 35062 40774 35076 40826
rect 35100 40774 35114 40826
rect 35114 40774 35126 40826
rect 35126 40774 35156 40826
rect 35180 40774 35190 40826
rect 35190 40774 35236 40826
rect 34940 40772 34996 40774
rect 35020 40772 35076 40774
rect 35100 40772 35156 40774
rect 35180 40772 35236 40774
rect 19580 40282 19636 40284
rect 19660 40282 19716 40284
rect 19740 40282 19796 40284
rect 19820 40282 19876 40284
rect 19580 40230 19626 40282
rect 19626 40230 19636 40282
rect 19660 40230 19690 40282
rect 19690 40230 19702 40282
rect 19702 40230 19716 40282
rect 19740 40230 19754 40282
rect 19754 40230 19766 40282
rect 19766 40230 19796 40282
rect 19820 40230 19830 40282
rect 19830 40230 19876 40282
rect 19580 40228 19636 40230
rect 19660 40228 19716 40230
rect 19740 40228 19796 40230
rect 19820 40228 19876 40230
rect 34940 39738 34996 39740
rect 35020 39738 35076 39740
rect 35100 39738 35156 39740
rect 35180 39738 35236 39740
rect 34940 39686 34986 39738
rect 34986 39686 34996 39738
rect 35020 39686 35050 39738
rect 35050 39686 35062 39738
rect 35062 39686 35076 39738
rect 35100 39686 35114 39738
rect 35114 39686 35126 39738
rect 35126 39686 35156 39738
rect 35180 39686 35190 39738
rect 35190 39686 35236 39738
rect 34940 39684 34996 39686
rect 35020 39684 35076 39686
rect 35100 39684 35156 39686
rect 35180 39684 35236 39686
rect 19580 39194 19636 39196
rect 19660 39194 19716 39196
rect 19740 39194 19796 39196
rect 19820 39194 19876 39196
rect 19580 39142 19626 39194
rect 19626 39142 19636 39194
rect 19660 39142 19690 39194
rect 19690 39142 19702 39194
rect 19702 39142 19716 39194
rect 19740 39142 19754 39194
rect 19754 39142 19766 39194
rect 19766 39142 19796 39194
rect 19820 39142 19830 39194
rect 19830 39142 19876 39194
rect 19580 39140 19636 39142
rect 19660 39140 19716 39142
rect 19740 39140 19796 39142
rect 19820 39140 19876 39142
rect 34940 38650 34996 38652
rect 35020 38650 35076 38652
rect 35100 38650 35156 38652
rect 35180 38650 35236 38652
rect 34940 38598 34986 38650
rect 34986 38598 34996 38650
rect 35020 38598 35050 38650
rect 35050 38598 35062 38650
rect 35062 38598 35076 38650
rect 35100 38598 35114 38650
rect 35114 38598 35126 38650
rect 35126 38598 35156 38650
rect 35180 38598 35190 38650
rect 35190 38598 35236 38650
rect 34940 38596 34996 38598
rect 35020 38596 35076 38598
rect 35100 38596 35156 38598
rect 35180 38596 35236 38598
rect 19580 38106 19636 38108
rect 19660 38106 19716 38108
rect 19740 38106 19796 38108
rect 19820 38106 19876 38108
rect 19580 38054 19626 38106
rect 19626 38054 19636 38106
rect 19660 38054 19690 38106
rect 19690 38054 19702 38106
rect 19702 38054 19716 38106
rect 19740 38054 19754 38106
rect 19754 38054 19766 38106
rect 19766 38054 19796 38106
rect 19820 38054 19830 38106
rect 19830 38054 19876 38106
rect 19580 38052 19636 38054
rect 19660 38052 19716 38054
rect 19740 38052 19796 38054
rect 19820 38052 19876 38054
rect 34940 37562 34996 37564
rect 35020 37562 35076 37564
rect 35100 37562 35156 37564
rect 35180 37562 35236 37564
rect 34940 37510 34986 37562
rect 34986 37510 34996 37562
rect 35020 37510 35050 37562
rect 35050 37510 35062 37562
rect 35062 37510 35076 37562
rect 35100 37510 35114 37562
rect 35114 37510 35126 37562
rect 35126 37510 35156 37562
rect 35180 37510 35190 37562
rect 35190 37510 35236 37562
rect 34940 37508 34996 37510
rect 35020 37508 35076 37510
rect 35100 37508 35156 37510
rect 35180 37508 35236 37510
rect 19580 37018 19636 37020
rect 19660 37018 19716 37020
rect 19740 37018 19796 37020
rect 19820 37018 19876 37020
rect 19580 36966 19626 37018
rect 19626 36966 19636 37018
rect 19660 36966 19690 37018
rect 19690 36966 19702 37018
rect 19702 36966 19716 37018
rect 19740 36966 19754 37018
rect 19754 36966 19766 37018
rect 19766 36966 19796 37018
rect 19820 36966 19830 37018
rect 19830 36966 19876 37018
rect 19580 36964 19636 36966
rect 19660 36964 19716 36966
rect 19740 36964 19796 36966
rect 19820 36964 19876 36966
rect 34940 36474 34996 36476
rect 35020 36474 35076 36476
rect 35100 36474 35156 36476
rect 35180 36474 35236 36476
rect 34940 36422 34986 36474
rect 34986 36422 34996 36474
rect 35020 36422 35050 36474
rect 35050 36422 35062 36474
rect 35062 36422 35076 36474
rect 35100 36422 35114 36474
rect 35114 36422 35126 36474
rect 35126 36422 35156 36474
rect 35180 36422 35190 36474
rect 35190 36422 35236 36474
rect 34940 36420 34996 36422
rect 35020 36420 35076 36422
rect 35100 36420 35156 36422
rect 35180 36420 35236 36422
rect 19580 35930 19636 35932
rect 19660 35930 19716 35932
rect 19740 35930 19796 35932
rect 19820 35930 19876 35932
rect 19580 35878 19626 35930
rect 19626 35878 19636 35930
rect 19660 35878 19690 35930
rect 19690 35878 19702 35930
rect 19702 35878 19716 35930
rect 19740 35878 19754 35930
rect 19754 35878 19766 35930
rect 19766 35878 19796 35930
rect 19820 35878 19830 35930
rect 19830 35878 19876 35930
rect 19580 35876 19636 35878
rect 19660 35876 19716 35878
rect 19740 35876 19796 35878
rect 19820 35876 19876 35878
rect 34940 35386 34996 35388
rect 35020 35386 35076 35388
rect 35100 35386 35156 35388
rect 35180 35386 35236 35388
rect 34940 35334 34986 35386
rect 34986 35334 34996 35386
rect 35020 35334 35050 35386
rect 35050 35334 35062 35386
rect 35062 35334 35076 35386
rect 35100 35334 35114 35386
rect 35114 35334 35126 35386
rect 35126 35334 35156 35386
rect 35180 35334 35190 35386
rect 35190 35334 35236 35386
rect 34940 35332 34996 35334
rect 35020 35332 35076 35334
rect 35100 35332 35156 35334
rect 35180 35332 35236 35334
rect 19580 34842 19636 34844
rect 19660 34842 19716 34844
rect 19740 34842 19796 34844
rect 19820 34842 19876 34844
rect 19580 34790 19626 34842
rect 19626 34790 19636 34842
rect 19660 34790 19690 34842
rect 19690 34790 19702 34842
rect 19702 34790 19716 34842
rect 19740 34790 19754 34842
rect 19754 34790 19766 34842
rect 19766 34790 19796 34842
rect 19820 34790 19830 34842
rect 19830 34790 19876 34842
rect 19580 34788 19636 34790
rect 19660 34788 19716 34790
rect 19740 34788 19796 34790
rect 19820 34788 19876 34790
rect 34940 34298 34996 34300
rect 35020 34298 35076 34300
rect 35100 34298 35156 34300
rect 35180 34298 35236 34300
rect 34940 34246 34986 34298
rect 34986 34246 34996 34298
rect 35020 34246 35050 34298
rect 35050 34246 35062 34298
rect 35062 34246 35076 34298
rect 35100 34246 35114 34298
rect 35114 34246 35126 34298
rect 35126 34246 35156 34298
rect 35180 34246 35190 34298
rect 35190 34246 35236 34298
rect 34940 34244 34996 34246
rect 35020 34244 35076 34246
rect 35100 34244 35156 34246
rect 35180 34244 35236 34246
rect 19580 33754 19636 33756
rect 19660 33754 19716 33756
rect 19740 33754 19796 33756
rect 19820 33754 19876 33756
rect 19580 33702 19626 33754
rect 19626 33702 19636 33754
rect 19660 33702 19690 33754
rect 19690 33702 19702 33754
rect 19702 33702 19716 33754
rect 19740 33702 19754 33754
rect 19754 33702 19766 33754
rect 19766 33702 19796 33754
rect 19820 33702 19830 33754
rect 19830 33702 19876 33754
rect 19580 33700 19636 33702
rect 19660 33700 19716 33702
rect 19740 33700 19796 33702
rect 19820 33700 19876 33702
rect 34940 33210 34996 33212
rect 35020 33210 35076 33212
rect 35100 33210 35156 33212
rect 35180 33210 35236 33212
rect 34940 33158 34986 33210
rect 34986 33158 34996 33210
rect 35020 33158 35050 33210
rect 35050 33158 35062 33210
rect 35062 33158 35076 33210
rect 35100 33158 35114 33210
rect 35114 33158 35126 33210
rect 35126 33158 35156 33210
rect 35180 33158 35190 33210
rect 35190 33158 35236 33210
rect 34940 33156 34996 33158
rect 35020 33156 35076 33158
rect 35100 33156 35156 33158
rect 35180 33156 35236 33158
rect 19580 32666 19636 32668
rect 19660 32666 19716 32668
rect 19740 32666 19796 32668
rect 19820 32666 19876 32668
rect 19580 32614 19626 32666
rect 19626 32614 19636 32666
rect 19660 32614 19690 32666
rect 19690 32614 19702 32666
rect 19702 32614 19716 32666
rect 19740 32614 19754 32666
rect 19754 32614 19766 32666
rect 19766 32614 19796 32666
rect 19820 32614 19830 32666
rect 19830 32614 19876 32666
rect 19580 32612 19636 32614
rect 19660 32612 19716 32614
rect 19740 32612 19796 32614
rect 19820 32612 19876 32614
rect 34940 32122 34996 32124
rect 35020 32122 35076 32124
rect 35100 32122 35156 32124
rect 35180 32122 35236 32124
rect 34940 32070 34986 32122
rect 34986 32070 34996 32122
rect 35020 32070 35050 32122
rect 35050 32070 35062 32122
rect 35062 32070 35076 32122
rect 35100 32070 35114 32122
rect 35114 32070 35126 32122
rect 35126 32070 35156 32122
rect 35180 32070 35190 32122
rect 35190 32070 35236 32122
rect 34940 32068 34996 32070
rect 35020 32068 35076 32070
rect 35100 32068 35156 32070
rect 35180 32068 35236 32070
rect 19580 31578 19636 31580
rect 19660 31578 19716 31580
rect 19740 31578 19796 31580
rect 19820 31578 19876 31580
rect 19580 31526 19626 31578
rect 19626 31526 19636 31578
rect 19660 31526 19690 31578
rect 19690 31526 19702 31578
rect 19702 31526 19716 31578
rect 19740 31526 19754 31578
rect 19754 31526 19766 31578
rect 19766 31526 19796 31578
rect 19820 31526 19830 31578
rect 19830 31526 19876 31578
rect 19580 31524 19636 31526
rect 19660 31524 19716 31526
rect 19740 31524 19796 31526
rect 19820 31524 19876 31526
rect 34940 31034 34996 31036
rect 35020 31034 35076 31036
rect 35100 31034 35156 31036
rect 35180 31034 35236 31036
rect 34940 30982 34986 31034
rect 34986 30982 34996 31034
rect 35020 30982 35050 31034
rect 35050 30982 35062 31034
rect 35062 30982 35076 31034
rect 35100 30982 35114 31034
rect 35114 30982 35126 31034
rect 35126 30982 35156 31034
rect 35180 30982 35190 31034
rect 35190 30982 35236 31034
rect 34940 30980 34996 30982
rect 35020 30980 35076 30982
rect 35100 30980 35156 30982
rect 35180 30980 35236 30982
rect 19580 30490 19636 30492
rect 19660 30490 19716 30492
rect 19740 30490 19796 30492
rect 19820 30490 19876 30492
rect 19580 30438 19626 30490
rect 19626 30438 19636 30490
rect 19660 30438 19690 30490
rect 19690 30438 19702 30490
rect 19702 30438 19716 30490
rect 19740 30438 19754 30490
rect 19754 30438 19766 30490
rect 19766 30438 19796 30490
rect 19820 30438 19830 30490
rect 19830 30438 19876 30490
rect 19580 30436 19636 30438
rect 19660 30436 19716 30438
rect 19740 30436 19796 30438
rect 19820 30436 19876 30438
rect 34940 29946 34996 29948
rect 35020 29946 35076 29948
rect 35100 29946 35156 29948
rect 35180 29946 35236 29948
rect 34940 29894 34986 29946
rect 34986 29894 34996 29946
rect 35020 29894 35050 29946
rect 35050 29894 35062 29946
rect 35062 29894 35076 29946
rect 35100 29894 35114 29946
rect 35114 29894 35126 29946
rect 35126 29894 35156 29946
rect 35180 29894 35190 29946
rect 35190 29894 35236 29946
rect 34940 29892 34996 29894
rect 35020 29892 35076 29894
rect 35100 29892 35156 29894
rect 35180 29892 35236 29894
rect 19580 29402 19636 29404
rect 19660 29402 19716 29404
rect 19740 29402 19796 29404
rect 19820 29402 19876 29404
rect 19580 29350 19626 29402
rect 19626 29350 19636 29402
rect 19660 29350 19690 29402
rect 19690 29350 19702 29402
rect 19702 29350 19716 29402
rect 19740 29350 19754 29402
rect 19754 29350 19766 29402
rect 19766 29350 19796 29402
rect 19820 29350 19830 29402
rect 19830 29350 19876 29402
rect 19580 29348 19636 29350
rect 19660 29348 19716 29350
rect 19740 29348 19796 29350
rect 19820 29348 19876 29350
rect 34940 28858 34996 28860
rect 35020 28858 35076 28860
rect 35100 28858 35156 28860
rect 35180 28858 35236 28860
rect 34940 28806 34986 28858
rect 34986 28806 34996 28858
rect 35020 28806 35050 28858
rect 35050 28806 35062 28858
rect 35062 28806 35076 28858
rect 35100 28806 35114 28858
rect 35114 28806 35126 28858
rect 35126 28806 35156 28858
rect 35180 28806 35190 28858
rect 35190 28806 35236 28858
rect 34940 28804 34996 28806
rect 35020 28804 35076 28806
rect 35100 28804 35156 28806
rect 35180 28804 35236 28806
rect 19580 28314 19636 28316
rect 19660 28314 19716 28316
rect 19740 28314 19796 28316
rect 19820 28314 19876 28316
rect 19580 28262 19626 28314
rect 19626 28262 19636 28314
rect 19660 28262 19690 28314
rect 19690 28262 19702 28314
rect 19702 28262 19716 28314
rect 19740 28262 19754 28314
rect 19754 28262 19766 28314
rect 19766 28262 19796 28314
rect 19820 28262 19830 28314
rect 19830 28262 19876 28314
rect 19580 28260 19636 28262
rect 19660 28260 19716 28262
rect 19740 28260 19796 28262
rect 19820 28260 19876 28262
rect 34940 27770 34996 27772
rect 35020 27770 35076 27772
rect 35100 27770 35156 27772
rect 35180 27770 35236 27772
rect 34940 27718 34986 27770
rect 34986 27718 34996 27770
rect 35020 27718 35050 27770
rect 35050 27718 35062 27770
rect 35062 27718 35076 27770
rect 35100 27718 35114 27770
rect 35114 27718 35126 27770
rect 35126 27718 35156 27770
rect 35180 27718 35190 27770
rect 35190 27718 35236 27770
rect 34940 27716 34996 27718
rect 35020 27716 35076 27718
rect 35100 27716 35156 27718
rect 35180 27716 35236 27718
rect 19580 27226 19636 27228
rect 19660 27226 19716 27228
rect 19740 27226 19796 27228
rect 19820 27226 19876 27228
rect 19580 27174 19626 27226
rect 19626 27174 19636 27226
rect 19660 27174 19690 27226
rect 19690 27174 19702 27226
rect 19702 27174 19716 27226
rect 19740 27174 19754 27226
rect 19754 27174 19766 27226
rect 19766 27174 19796 27226
rect 19820 27174 19830 27226
rect 19830 27174 19876 27226
rect 19580 27172 19636 27174
rect 19660 27172 19716 27174
rect 19740 27172 19796 27174
rect 19820 27172 19876 27174
rect 34940 26682 34996 26684
rect 35020 26682 35076 26684
rect 35100 26682 35156 26684
rect 35180 26682 35236 26684
rect 34940 26630 34986 26682
rect 34986 26630 34996 26682
rect 35020 26630 35050 26682
rect 35050 26630 35062 26682
rect 35062 26630 35076 26682
rect 35100 26630 35114 26682
rect 35114 26630 35126 26682
rect 35126 26630 35156 26682
rect 35180 26630 35190 26682
rect 35190 26630 35236 26682
rect 34940 26628 34996 26630
rect 35020 26628 35076 26630
rect 35100 26628 35156 26630
rect 35180 26628 35236 26630
rect 19580 26138 19636 26140
rect 19660 26138 19716 26140
rect 19740 26138 19796 26140
rect 19820 26138 19876 26140
rect 19580 26086 19626 26138
rect 19626 26086 19636 26138
rect 19660 26086 19690 26138
rect 19690 26086 19702 26138
rect 19702 26086 19716 26138
rect 19740 26086 19754 26138
rect 19754 26086 19766 26138
rect 19766 26086 19796 26138
rect 19820 26086 19830 26138
rect 19830 26086 19876 26138
rect 19580 26084 19636 26086
rect 19660 26084 19716 26086
rect 19740 26084 19796 26086
rect 19820 26084 19876 26086
rect 34940 25594 34996 25596
rect 35020 25594 35076 25596
rect 35100 25594 35156 25596
rect 35180 25594 35236 25596
rect 34940 25542 34986 25594
rect 34986 25542 34996 25594
rect 35020 25542 35050 25594
rect 35050 25542 35062 25594
rect 35062 25542 35076 25594
rect 35100 25542 35114 25594
rect 35114 25542 35126 25594
rect 35126 25542 35156 25594
rect 35180 25542 35190 25594
rect 35190 25542 35236 25594
rect 34940 25540 34996 25542
rect 35020 25540 35076 25542
rect 35100 25540 35156 25542
rect 35180 25540 35236 25542
rect 19580 25050 19636 25052
rect 19660 25050 19716 25052
rect 19740 25050 19796 25052
rect 19820 25050 19876 25052
rect 19580 24998 19626 25050
rect 19626 24998 19636 25050
rect 19660 24998 19690 25050
rect 19690 24998 19702 25050
rect 19702 24998 19716 25050
rect 19740 24998 19754 25050
rect 19754 24998 19766 25050
rect 19766 24998 19796 25050
rect 19820 24998 19830 25050
rect 19830 24998 19876 25050
rect 19580 24996 19636 24998
rect 19660 24996 19716 24998
rect 19740 24996 19796 24998
rect 19820 24996 19876 24998
rect 34940 24506 34996 24508
rect 35020 24506 35076 24508
rect 35100 24506 35156 24508
rect 35180 24506 35236 24508
rect 34940 24454 34986 24506
rect 34986 24454 34996 24506
rect 35020 24454 35050 24506
rect 35050 24454 35062 24506
rect 35062 24454 35076 24506
rect 35100 24454 35114 24506
rect 35114 24454 35126 24506
rect 35126 24454 35156 24506
rect 35180 24454 35190 24506
rect 35190 24454 35236 24506
rect 34940 24452 34996 24454
rect 35020 24452 35076 24454
rect 35100 24452 35156 24454
rect 35180 24452 35236 24454
rect 19580 23962 19636 23964
rect 19660 23962 19716 23964
rect 19740 23962 19796 23964
rect 19820 23962 19876 23964
rect 19580 23910 19626 23962
rect 19626 23910 19636 23962
rect 19660 23910 19690 23962
rect 19690 23910 19702 23962
rect 19702 23910 19716 23962
rect 19740 23910 19754 23962
rect 19754 23910 19766 23962
rect 19766 23910 19796 23962
rect 19820 23910 19830 23962
rect 19830 23910 19876 23962
rect 19580 23908 19636 23910
rect 19660 23908 19716 23910
rect 19740 23908 19796 23910
rect 19820 23908 19876 23910
rect 34940 23418 34996 23420
rect 35020 23418 35076 23420
rect 35100 23418 35156 23420
rect 35180 23418 35236 23420
rect 34940 23366 34986 23418
rect 34986 23366 34996 23418
rect 35020 23366 35050 23418
rect 35050 23366 35062 23418
rect 35062 23366 35076 23418
rect 35100 23366 35114 23418
rect 35114 23366 35126 23418
rect 35126 23366 35156 23418
rect 35180 23366 35190 23418
rect 35190 23366 35236 23418
rect 34940 23364 34996 23366
rect 35020 23364 35076 23366
rect 35100 23364 35156 23366
rect 35180 23364 35236 23366
rect 19580 22874 19636 22876
rect 19660 22874 19716 22876
rect 19740 22874 19796 22876
rect 19820 22874 19876 22876
rect 19580 22822 19626 22874
rect 19626 22822 19636 22874
rect 19660 22822 19690 22874
rect 19690 22822 19702 22874
rect 19702 22822 19716 22874
rect 19740 22822 19754 22874
rect 19754 22822 19766 22874
rect 19766 22822 19796 22874
rect 19820 22822 19830 22874
rect 19830 22822 19876 22874
rect 19580 22820 19636 22822
rect 19660 22820 19716 22822
rect 19740 22820 19796 22822
rect 19820 22820 19876 22822
rect 34940 22330 34996 22332
rect 35020 22330 35076 22332
rect 35100 22330 35156 22332
rect 35180 22330 35236 22332
rect 34940 22278 34986 22330
rect 34986 22278 34996 22330
rect 35020 22278 35050 22330
rect 35050 22278 35062 22330
rect 35062 22278 35076 22330
rect 35100 22278 35114 22330
rect 35114 22278 35126 22330
rect 35126 22278 35156 22330
rect 35180 22278 35190 22330
rect 35190 22278 35236 22330
rect 34940 22276 34996 22278
rect 35020 22276 35076 22278
rect 35100 22276 35156 22278
rect 35180 22276 35236 22278
rect 19580 21786 19636 21788
rect 19660 21786 19716 21788
rect 19740 21786 19796 21788
rect 19820 21786 19876 21788
rect 19580 21734 19626 21786
rect 19626 21734 19636 21786
rect 19660 21734 19690 21786
rect 19690 21734 19702 21786
rect 19702 21734 19716 21786
rect 19740 21734 19754 21786
rect 19754 21734 19766 21786
rect 19766 21734 19796 21786
rect 19820 21734 19830 21786
rect 19830 21734 19876 21786
rect 19580 21732 19636 21734
rect 19660 21732 19716 21734
rect 19740 21732 19796 21734
rect 19820 21732 19876 21734
rect 34940 21242 34996 21244
rect 35020 21242 35076 21244
rect 35100 21242 35156 21244
rect 35180 21242 35236 21244
rect 34940 21190 34986 21242
rect 34986 21190 34996 21242
rect 35020 21190 35050 21242
rect 35050 21190 35062 21242
rect 35062 21190 35076 21242
rect 35100 21190 35114 21242
rect 35114 21190 35126 21242
rect 35126 21190 35156 21242
rect 35180 21190 35190 21242
rect 35190 21190 35236 21242
rect 34940 21188 34996 21190
rect 35020 21188 35076 21190
rect 35100 21188 35156 21190
rect 35180 21188 35236 21190
rect 19580 20698 19636 20700
rect 19660 20698 19716 20700
rect 19740 20698 19796 20700
rect 19820 20698 19876 20700
rect 19580 20646 19626 20698
rect 19626 20646 19636 20698
rect 19660 20646 19690 20698
rect 19690 20646 19702 20698
rect 19702 20646 19716 20698
rect 19740 20646 19754 20698
rect 19754 20646 19766 20698
rect 19766 20646 19796 20698
rect 19820 20646 19830 20698
rect 19830 20646 19876 20698
rect 19580 20644 19636 20646
rect 19660 20644 19716 20646
rect 19740 20644 19796 20646
rect 19820 20644 19876 20646
rect 34940 20154 34996 20156
rect 35020 20154 35076 20156
rect 35100 20154 35156 20156
rect 35180 20154 35236 20156
rect 34940 20102 34986 20154
rect 34986 20102 34996 20154
rect 35020 20102 35050 20154
rect 35050 20102 35062 20154
rect 35062 20102 35076 20154
rect 35100 20102 35114 20154
rect 35114 20102 35126 20154
rect 35126 20102 35156 20154
rect 35180 20102 35190 20154
rect 35190 20102 35236 20154
rect 34940 20100 34996 20102
rect 35020 20100 35076 20102
rect 35100 20100 35156 20102
rect 35180 20100 35236 20102
rect 19580 19610 19636 19612
rect 19660 19610 19716 19612
rect 19740 19610 19796 19612
rect 19820 19610 19876 19612
rect 19580 19558 19626 19610
rect 19626 19558 19636 19610
rect 19660 19558 19690 19610
rect 19690 19558 19702 19610
rect 19702 19558 19716 19610
rect 19740 19558 19754 19610
rect 19754 19558 19766 19610
rect 19766 19558 19796 19610
rect 19820 19558 19830 19610
rect 19830 19558 19876 19610
rect 19580 19556 19636 19558
rect 19660 19556 19716 19558
rect 19740 19556 19796 19558
rect 19820 19556 19876 19558
rect 34940 19066 34996 19068
rect 35020 19066 35076 19068
rect 35100 19066 35156 19068
rect 35180 19066 35236 19068
rect 34940 19014 34986 19066
rect 34986 19014 34996 19066
rect 35020 19014 35050 19066
rect 35050 19014 35062 19066
rect 35062 19014 35076 19066
rect 35100 19014 35114 19066
rect 35114 19014 35126 19066
rect 35126 19014 35156 19066
rect 35180 19014 35190 19066
rect 35190 19014 35236 19066
rect 34940 19012 34996 19014
rect 35020 19012 35076 19014
rect 35100 19012 35156 19014
rect 35180 19012 35236 19014
rect 19580 18522 19636 18524
rect 19660 18522 19716 18524
rect 19740 18522 19796 18524
rect 19820 18522 19876 18524
rect 19580 18470 19626 18522
rect 19626 18470 19636 18522
rect 19660 18470 19690 18522
rect 19690 18470 19702 18522
rect 19702 18470 19716 18522
rect 19740 18470 19754 18522
rect 19754 18470 19766 18522
rect 19766 18470 19796 18522
rect 19820 18470 19830 18522
rect 19830 18470 19876 18522
rect 19580 18468 19636 18470
rect 19660 18468 19716 18470
rect 19740 18468 19796 18470
rect 19820 18468 19876 18470
rect 34940 17978 34996 17980
rect 35020 17978 35076 17980
rect 35100 17978 35156 17980
rect 35180 17978 35236 17980
rect 34940 17926 34986 17978
rect 34986 17926 34996 17978
rect 35020 17926 35050 17978
rect 35050 17926 35062 17978
rect 35062 17926 35076 17978
rect 35100 17926 35114 17978
rect 35114 17926 35126 17978
rect 35126 17926 35156 17978
rect 35180 17926 35190 17978
rect 35190 17926 35236 17978
rect 34940 17924 34996 17926
rect 35020 17924 35076 17926
rect 35100 17924 35156 17926
rect 35180 17924 35236 17926
rect 19580 17434 19636 17436
rect 19660 17434 19716 17436
rect 19740 17434 19796 17436
rect 19820 17434 19876 17436
rect 19580 17382 19626 17434
rect 19626 17382 19636 17434
rect 19660 17382 19690 17434
rect 19690 17382 19702 17434
rect 19702 17382 19716 17434
rect 19740 17382 19754 17434
rect 19754 17382 19766 17434
rect 19766 17382 19796 17434
rect 19820 17382 19830 17434
rect 19830 17382 19876 17434
rect 19580 17380 19636 17382
rect 19660 17380 19716 17382
rect 19740 17380 19796 17382
rect 19820 17380 19876 17382
rect 34940 16890 34996 16892
rect 35020 16890 35076 16892
rect 35100 16890 35156 16892
rect 35180 16890 35236 16892
rect 34940 16838 34986 16890
rect 34986 16838 34996 16890
rect 35020 16838 35050 16890
rect 35050 16838 35062 16890
rect 35062 16838 35076 16890
rect 35100 16838 35114 16890
rect 35114 16838 35126 16890
rect 35126 16838 35156 16890
rect 35180 16838 35190 16890
rect 35190 16838 35236 16890
rect 34940 16836 34996 16838
rect 35020 16836 35076 16838
rect 35100 16836 35156 16838
rect 35180 16836 35236 16838
rect 19580 16346 19636 16348
rect 19660 16346 19716 16348
rect 19740 16346 19796 16348
rect 19820 16346 19876 16348
rect 19580 16294 19626 16346
rect 19626 16294 19636 16346
rect 19660 16294 19690 16346
rect 19690 16294 19702 16346
rect 19702 16294 19716 16346
rect 19740 16294 19754 16346
rect 19754 16294 19766 16346
rect 19766 16294 19796 16346
rect 19820 16294 19830 16346
rect 19830 16294 19876 16346
rect 19580 16292 19636 16294
rect 19660 16292 19716 16294
rect 19740 16292 19796 16294
rect 19820 16292 19876 16294
rect 34940 15802 34996 15804
rect 35020 15802 35076 15804
rect 35100 15802 35156 15804
rect 35180 15802 35236 15804
rect 34940 15750 34986 15802
rect 34986 15750 34996 15802
rect 35020 15750 35050 15802
rect 35050 15750 35062 15802
rect 35062 15750 35076 15802
rect 35100 15750 35114 15802
rect 35114 15750 35126 15802
rect 35126 15750 35156 15802
rect 35180 15750 35190 15802
rect 35190 15750 35236 15802
rect 34940 15748 34996 15750
rect 35020 15748 35076 15750
rect 35100 15748 35156 15750
rect 35180 15748 35236 15750
rect 19580 15258 19636 15260
rect 19660 15258 19716 15260
rect 19740 15258 19796 15260
rect 19820 15258 19876 15260
rect 19580 15206 19626 15258
rect 19626 15206 19636 15258
rect 19660 15206 19690 15258
rect 19690 15206 19702 15258
rect 19702 15206 19716 15258
rect 19740 15206 19754 15258
rect 19754 15206 19766 15258
rect 19766 15206 19796 15258
rect 19820 15206 19830 15258
rect 19830 15206 19876 15258
rect 19580 15204 19636 15206
rect 19660 15204 19716 15206
rect 19740 15204 19796 15206
rect 19820 15204 19876 15206
rect 34940 14714 34996 14716
rect 35020 14714 35076 14716
rect 35100 14714 35156 14716
rect 35180 14714 35236 14716
rect 34940 14662 34986 14714
rect 34986 14662 34996 14714
rect 35020 14662 35050 14714
rect 35050 14662 35062 14714
rect 35062 14662 35076 14714
rect 35100 14662 35114 14714
rect 35114 14662 35126 14714
rect 35126 14662 35156 14714
rect 35180 14662 35190 14714
rect 35190 14662 35236 14714
rect 34940 14660 34996 14662
rect 35020 14660 35076 14662
rect 35100 14660 35156 14662
rect 35180 14660 35236 14662
rect 19580 14170 19636 14172
rect 19660 14170 19716 14172
rect 19740 14170 19796 14172
rect 19820 14170 19876 14172
rect 19580 14118 19626 14170
rect 19626 14118 19636 14170
rect 19660 14118 19690 14170
rect 19690 14118 19702 14170
rect 19702 14118 19716 14170
rect 19740 14118 19754 14170
rect 19754 14118 19766 14170
rect 19766 14118 19796 14170
rect 19820 14118 19830 14170
rect 19830 14118 19876 14170
rect 19580 14116 19636 14118
rect 19660 14116 19716 14118
rect 19740 14116 19796 14118
rect 19820 14116 19876 14118
rect 34940 13626 34996 13628
rect 35020 13626 35076 13628
rect 35100 13626 35156 13628
rect 35180 13626 35236 13628
rect 34940 13574 34986 13626
rect 34986 13574 34996 13626
rect 35020 13574 35050 13626
rect 35050 13574 35062 13626
rect 35062 13574 35076 13626
rect 35100 13574 35114 13626
rect 35114 13574 35126 13626
rect 35126 13574 35156 13626
rect 35180 13574 35190 13626
rect 35190 13574 35236 13626
rect 34940 13572 34996 13574
rect 35020 13572 35076 13574
rect 35100 13572 35156 13574
rect 35180 13572 35236 13574
rect 19580 13082 19636 13084
rect 19660 13082 19716 13084
rect 19740 13082 19796 13084
rect 19820 13082 19876 13084
rect 19580 13030 19626 13082
rect 19626 13030 19636 13082
rect 19660 13030 19690 13082
rect 19690 13030 19702 13082
rect 19702 13030 19716 13082
rect 19740 13030 19754 13082
rect 19754 13030 19766 13082
rect 19766 13030 19796 13082
rect 19820 13030 19830 13082
rect 19830 13030 19876 13082
rect 19580 13028 19636 13030
rect 19660 13028 19716 13030
rect 19740 13028 19796 13030
rect 19820 13028 19876 13030
rect 34940 12538 34996 12540
rect 35020 12538 35076 12540
rect 35100 12538 35156 12540
rect 35180 12538 35236 12540
rect 34940 12486 34986 12538
rect 34986 12486 34996 12538
rect 35020 12486 35050 12538
rect 35050 12486 35062 12538
rect 35062 12486 35076 12538
rect 35100 12486 35114 12538
rect 35114 12486 35126 12538
rect 35126 12486 35156 12538
rect 35180 12486 35190 12538
rect 35190 12486 35236 12538
rect 34940 12484 34996 12486
rect 35020 12484 35076 12486
rect 35100 12484 35156 12486
rect 35180 12484 35236 12486
rect 19580 11994 19636 11996
rect 19660 11994 19716 11996
rect 19740 11994 19796 11996
rect 19820 11994 19876 11996
rect 19580 11942 19626 11994
rect 19626 11942 19636 11994
rect 19660 11942 19690 11994
rect 19690 11942 19702 11994
rect 19702 11942 19716 11994
rect 19740 11942 19754 11994
rect 19754 11942 19766 11994
rect 19766 11942 19796 11994
rect 19820 11942 19830 11994
rect 19830 11942 19876 11994
rect 19580 11940 19636 11942
rect 19660 11940 19716 11942
rect 19740 11940 19796 11942
rect 19820 11940 19876 11942
rect 34940 11450 34996 11452
rect 35020 11450 35076 11452
rect 35100 11450 35156 11452
rect 35180 11450 35236 11452
rect 34940 11398 34986 11450
rect 34986 11398 34996 11450
rect 35020 11398 35050 11450
rect 35050 11398 35062 11450
rect 35062 11398 35076 11450
rect 35100 11398 35114 11450
rect 35114 11398 35126 11450
rect 35126 11398 35156 11450
rect 35180 11398 35190 11450
rect 35190 11398 35236 11450
rect 34940 11396 34996 11398
rect 35020 11396 35076 11398
rect 35100 11396 35156 11398
rect 35180 11396 35236 11398
rect 19580 10906 19636 10908
rect 19660 10906 19716 10908
rect 19740 10906 19796 10908
rect 19820 10906 19876 10908
rect 19580 10854 19626 10906
rect 19626 10854 19636 10906
rect 19660 10854 19690 10906
rect 19690 10854 19702 10906
rect 19702 10854 19716 10906
rect 19740 10854 19754 10906
rect 19754 10854 19766 10906
rect 19766 10854 19796 10906
rect 19820 10854 19830 10906
rect 19830 10854 19876 10906
rect 19580 10852 19636 10854
rect 19660 10852 19716 10854
rect 19740 10852 19796 10854
rect 19820 10852 19876 10854
rect 34940 10362 34996 10364
rect 35020 10362 35076 10364
rect 35100 10362 35156 10364
rect 35180 10362 35236 10364
rect 34940 10310 34986 10362
rect 34986 10310 34996 10362
rect 35020 10310 35050 10362
rect 35050 10310 35062 10362
rect 35062 10310 35076 10362
rect 35100 10310 35114 10362
rect 35114 10310 35126 10362
rect 35126 10310 35156 10362
rect 35180 10310 35190 10362
rect 35190 10310 35236 10362
rect 34940 10308 34996 10310
rect 35020 10308 35076 10310
rect 35100 10308 35156 10310
rect 35180 10308 35236 10310
rect 19580 9818 19636 9820
rect 19660 9818 19716 9820
rect 19740 9818 19796 9820
rect 19820 9818 19876 9820
rect 19580 9766 19626 9818
rect 19626 9766 19636 9818
rect 19660 9766 19690 9818
rect 19690 9766 19702 9818
rect 19702 9766 19716 9818
rect 19740 9766 19754 9818
rect 19754 9766 19766 9818
rect 19766 9766 19796 9818
rect 19820 9766 19830 9818
rect 19830 9766 19876 9818
rect 19580 9764 19636 9766
rect 19660 9764 19716 9766
rect 19740 9764 19796 9766
rect 19820 9764 19876 9766
rect 34940 9274 34996 9276
rect 35020 9274 35076 9276
rect 35100 9274 35156 9276
rect 35180 9274 35236 9276
rect 34940 9222 34986 9274
rect 34986 9222 34996 9274
rect 35020 9222 35050 9274
rect 35050 9222 35062 9274
rect 35062 9222 35076 9274
rect 35100 9222 35114 9274
rect 35114 9222 35126 9274
rect 35126 9222 35156 9274
rect 35180 9222 35190 9274
rect 35190 9222 35236 9274
rect 34940 9220 34996 9222
rect 35020 9220 35076 9222
rect 35100 9220 35156 9222
rect 35180 9220 35236 9222
rect 19580 8730 19636 8732
rect 19660 8730 19716 8732
rect 19740 8730 19796 8732
rect 19820 8730 19876 8732
rect 19580 8678 19626 8730
rect 19626 8678 19636 8730
rect 19660 8678 19690 8730
rect 19690 8678 19702 8730
rect 19702 8678 19716 8730
rect 19740 8678 19754 8730
rect 19754 8678 19766 8730
rect 19766 8678 19796 8730
rect 19820 8678 19830 8730
rect 19830 8678 19876 8730
rect 19580 8676 19636 8678
rect 19660 8676 19716 8678
rect 19740 8676 19796 8678
rect 19820 8676 19876 8678
rect 34940 8186 34996 8188
rect 35020 8186 35076 8188
rect 35100 8186 35156 8188
rect 35180 8186 35236 8188
rect 34940 8134 34986 8186
rect 34986 8134 34996 8186
rect 35020 8134 35050 8186
rect 35050 8134 35062 8186
rect 35062 8134 35076 8186
rect 35100 8134 35114 8186
rect 35114 8134 35126 8186
rect 35126 8134 35156 8186
rect 35180 8134 35190 8186
rect 35190 8134 35236 8186
rect 34940 8132 34996 8134
rect 35020 8132 35076 8134
rect 35100 8132 35156 8134
rect 35180 8132 35236 8134
rect 19580 7642 19636 7644
rect 19660 7642 19716 7644
rect 19740 7642 19796 7644
rect 19820 7642 19876 7644
rect 19580 7590 19626 7642
rect 19626 7590 19636 7642
rect 19660 7590 19690 7642
rect 19690 7590 19702 7642
rect 19702 7590 19716 7642
rect 19740 7590 19754 7642
rect 19754 7590 19766 7642
rect 19766 7590 19796 7642
rect 19820 7590 19830 7642
rect 19830 7590 19876 7642
rect 19580 7588 19636 7590
rect 19660 7588 19716 7590
rect 19740 7588 19796 7590
rect 19820 7588 19876 7590
rect 34940 7098 34996 7100
rect 35020 7098 35076 7100
rect 35100 7098 35156 7100
rect 35180 7098 35236 7100
rect 34940 7046 34986 7098
rect 34986 7046 34996 7098
rect 35020 7046 35050 7098
rect 35050 7046 35062 7098
rect 35062 7046 35076 7098
rect 35100 7046 35114 7098
rect 35114 7046 35126 7098
rect 35126 7046 35156 7098
rect 35180 7046 35190 7098
rect 35190 7046 35236 7098
rect 34940 7044 34996 7046
rect 35020 7044 35076 7046
rect 35100 7044 35156 7046
rect 35180 7044 35236 7046
rect 19580 6554 19636 6556
rect 19660 6554 19716 6556
rect 19740 6554 19796 6556
rect 19820 6554 19876 6556
rect 19580 6502 19626 6554
rect 19626 6502 19636 6554
rect 19660 6502 19690 6554
rect 19690 6502 19702 6554
rect 19702 6502 19716 6554
rect 19740 6502 19754 6554
rect 19754 6502 19766 6554
rect 19766 6502 19796 6554
rect 19820 6502 19830 6554
rect 19830 6502 19876 6554
rect 19580 6500 19636 6502
rect 19660 6500 19716 6502
rect 19740 6500 19796 6502
rect 19820 6500 19876 6502
rect 34940 6010 34996 6012
rect 35020 6010 35076 6012
rect 35100 6010 35156 6012
rect 35180 6010 35236 6012
rect 34940 5958 34986 6010
rect 34986 5958 34996 6010
rect 35020 5958 35050 6010
rect 35050 5958 35062 6010
rect 35062 5958 35076 6010
rect 35100 5958 35114 6010
rect 35114 5958 35126 6010
rect 35126 5958 35156 6010
rect 35180 5958 35190 6010
rect 35190 5958 35236 6010
rect 34940 5956 34996 5958
rect 35020 5956 35076 5958
rect 35100 5956 35156 5958
rect 35180 5956 35236 5958
rect 19580 5466 19636 5468
rect 19660 5466 19716 5468
rect 19740 5466 19796 5468
rect 19820 5466 19876 5468
rect 19580 5414 19626 5466
rect 19626 5414 19636 5466
rect 19660 5414 19690 5466
rect 19690 5414 19702 5466
rect 19702 5414 19716 5466
rect 19740 5414 19754 5466
rect 19754 5414 19766 5466
rect 19766 5414 19796 5466
rect 19820 5414 19830 5466
rect 19830 5414 19876 5466
rect 19580 5412 19636 5414
rect 19660 5412 19716 5414
rect 19740 5412 19796 5414
rect 19820 5412 19876 5414
rect 34940 4922 34996 4924
rect 35020 4922 35076 4924
rect 35100 4922 35156 4924
rect 35180 4922 35236 4924
rect 34940 4870 34986 4922
rect 34986 4870 34996 4922
rect 35020 4870 35050 4922
rect 35050 4870 35062 4922
rect 35062 4870 35076 4922
rect 35100 4870 35114 4922
rect 35114 4870 35126 4922
rect 35126 4870 35156 4922
rect 35180 4870 35190 4922
rect 35190 4870 35236 4922
rect 34940 4868 34996 4870
rect 35020 4868 35076 4870
rect 35100 4868 35156 4870
rect 35180 4868 35236 4870
rect 4220 3834 4276 3836
rect 4300 3834 4356 3836
rect 4380 3834 4436 3836
rect 4460 3834 4516 3836
rect 4220 3782 4266 3834
rect 4266 3782 4276 3834
rect 4300 3782 4330 3834
rect 4330 3782 4342 3834
rect 4342 3782 4356 3834
rect 4380 3782 4394 3834
rect 4394 3782 4406 3834
rect 4406 3782 4436 3834
rect 4460 3782 4470 3834
rect 4470 3782 4516 3834
rect 4220 3780 4276 3782
rect 4300 3780 4356 3782
rect 4380 3780 4436 3782
rect 4460 3780 4516 3782
rect 4220 2746 4276 2748
rect 4300 2746 4356 2748
rect 4380 2746 4436 2748
rect 4460 2746 4516 2748
rect 4220 2694 4266 2746
rect 4266 2694 4276 2746
rect 4300 2694 4330 2746
rect 4330 2694 4342 2746
rect 4342 2694 4356 2746
rect 4380 2694 4394 2746
rect 4394 2694 4406 2746
rect 4406 2694 4436 2746
rect 4460 2694 4470 2746
rect 4470 2694 4516 2746
rect 4220 2692 4276 2694
rect 4300 2692 4356 2694
rect 4380 2692 4436 2694
rect 4460 2692 4516 2694
rect 19580 4378 19636 4380
rect 19660 4378 19716 4380
rect 19740 4378 19796 4380
rect 19820 4378 19876 4380
rect 19580 4326 19626 4378
rect 19626 4326 19636 4378
rect 19660 4326 19690 4378
rect 19690 4326 19702 4378
rect 19702 4326 19716 4378
rect 19740 4326 19754 4378
rect 19754 4326 19766 4378
rect 19766 4326 19796 4378
rect 19820 4326 19830 4378
rect 19830 4326 19876 4378
rect 19580 4324 19636 4326
rect 19660 4324 19716 4326
rect 19740 4324 19796 4326
rect 19820 4324 19876 4326
rect 34940 3834 34996 3836
rect 35020 3834 35076 3836
rect 35100 3834 35156 3836
rect 35180 3834 35236 3836
rect 34940 3782 34986 3834
rect 34986 3782 34996 3834
rect 35020 3782 35050 3834
rect 35050 3782 35062 3834
rect 35062 3782 35076 3834
rect 35100 3782 35114 3834
rect 35114 3782 35126 3834
rect 35126 3782 35156 3834
rect 35180 3782 35190 3834
rect 35190 3782 35236 3834
rect 34940 3780 34996 3782
rect 35020 3780 35076 3782
rect 35100 3780 35156 3782
rect 35180 3780 35236 3782
rect 19580 3290 19636 3292
rect 19660 3290 19716 3292
rect 19740 3290 19796 3292
rect 19820 3290 19876 3292
rect 19580 3238 19626 3290
rect 19626 3238 19636 3290
rect 19660 3238 19690 3290
rect 19690 3238 19702 3290
rect 19702 3238 19716 3290
rect 19740 3238 19754 3290
rect 19754 3238 19766 3290
rect 19766 3238 19796 3290
rect 19820 3238 19830 3290
rect 19830 3238 19876 3290
rect 19580 3236 19636 3238
rect 19660 3236 19716 3238
rect 19740 3236 19796 3238
rect 19820 3236 19876 3238
rect 19580 2202 19636 2204
rect 19660 2202 19716 2204
rect 19740 2202 19796 2204
rect 19820 2202 19876 2204
rect 19580 2150 19626 2202
rect 19626 2150 19636 2202
rect 19660 2150 19690 2202
rect 19690 2150 19702 2202
rect 19702 2150 19716 2202
rect 19740 2150 19754 2202
rect 19754 2150 19766 2202
rect 19766 2150 19796 2202
rect 19820 2150 19830 2202
rect 19830 2150 19876 2202
rect 19580 2148 19636 2150
rect 19660 2148 19716 2150
rect 19740 2148 19796 2150
rect 19820 2148 19876 2150
rect 34940 2746 34996 2748
rect 35020 2746 35076 2748
rect 35100 2746 35156 2748
rect 35180 2746 35236 2748
rect 34940 2694 34986 2746
rect 34986 2694 34996 2746
rect 35020 2694 35050 2746
rect 35050 2694 35062 2746
rect 35062 2694 35076 2746
rect 35100 2694 35114 2746
rect 35114 2694 35126 2746
rect 35126 2694 35156 2746
rect 35180 2694 35190 2746
rect 35190 2694 35236 2746
rect 34940 2692 34996 2694
rect 35020 2692 35076 2694
rect 35100 2692 35156 2694
rect 35180 2692 35236 2694
rect 50300 48986 50356 48988
rect 50380 48986 50436 48988
rect 50460 48986 50516 48988
rect 50540 48986 50596 48988
rect 50300 48934 50346 48986
rect 50346 48934 50356 48986
rect 50380 48934 50410 48986
rect 50410 48934 50422 48986
rect 50422 48934 50436 48986
rect 50460 48934 50474 48986
rect 50474 48934 50486 48986
rect 50486 48934 50516 48986
rect 50540 48934 50550 48986
rect 50550 48934 50596 48986
rect 50300 48932 50356 48934
rect 50380 48932 50436 48934
rect 50460 48932 50516 48934
rect 50540 48932 50596 48934
rect 50300 47898 50356 47900
rect 50380 47898 50436 47900
rect 50460 47898 50516 47900
rect 50540 47898 50596 47900
rect 50300 47846 50346 47898
rect 50346 47846 50356 47898
rect 50380 47846 50410 47898
rect 50410 47846 50422 47898
rect 50422 47846 50436 47898
rect 50460 47846 50474 47898
rect 50474 47846 50486 47898
rect 50486 47846 50516 47898
rect 50540 47846 50550 47898
rect 50550 47846 50596 47898
rect 50300 47844 50356 47846
rect 50380 47844 50436 47846
rect 50460 47844 50516 47846
rect 50540 47844 50596 47846
rect 50300 46810 50356 46812
rect 50380 46810 50436 46812
rect 50460 46810 50516 46812
rect 50540 46810 50596 46812
rect 50300 46758 50346 46810
rect 50346 46758 50356 46810
rect 50380 46758 50410 46810
rect 50410 46758 50422 46810
rect 50422 46758 50436 46810
rect 50460 46758 50474 46810
rect 50474 46758 50486 46810
rect 50486 46758 50516 46810
rect 50540 46758 50550 46810
rect 50550 46758 50596 46810
rect 50300 46756 50356 46758
rect 50380 46756 50436 46758
rect 50460 46756 50516 46758
rect 50540 46756 50596 46758
rect 50300 45722 50356 45724
rect 50380 45722 50436 45724
rect 50460 45722 50516 45724
rect 50540 45722 50596 45724
rect 50300 45670 50346 45722
rect 50346 45670 50356 45722
rect 50380 45670 50410 45722
rect 50410 45670 50422 45722
rect 50422 45670 50436 45722
rect 50460 45670 50474 45722
rect 50474 45670 50486 45722
rect 50486 45670 50516 45722
rect 50540 45670 50550 45722
rect 50550 45670 50596 45722
rect 50300 45668 50356 45670
rect 50380 45668 50436 45670
rect 50460 45668 50516 45670
rect 50540 45668 50596 45670
rect 50300 44634 50356 44636
rect 50380 44634 50436 44636
rect 50460 44634 50516 44636
rect 50540 44634 50596 44636
rect 50300 44582 50346 44634
rect 50346 44582 50356 44634
rect 50380 44582 50410 44634
rect 50410 44582 50422 44634
rect 50422 44582 50436 44634
rect 50460 44582 50474 44634
rect 50474 44582 50486 44634
rect 50486 44582 50516 44634
rect 50540 44582 50550 44634
rect 50550 44582 50596 44634
rect 50300 44580 50356 44582
rect 50380 44580 50436 44582
rect 50460 44580 50516 44582
rect 50540 44580 50596 44582
rect 50986 45464 51042 45520
rect 52642 45464 52698 45520
rect 50300 43546 50356 43548
rect 50380 43546 50436 43548
rect 50460 43546 50516 43548
rect 50540 43546 50596 43548
rect 50300 43494 50346 43546
rect 50346 43494 50356 43546
rect 50380 43494 50410 43546
rect 50410 43494 50422 43546
rect 50422 43494 50436 43546
rect 50460 43494 50474 43546
rect 50474 43494 50486 43546
rect 50486 43494 50516 43546
rect 50540 43494 50550 43546
rect 50550 43494 50596 43546
rect 50300 43492 50356 43494
rect 50380 43492 50436 43494
rect 50460 43492 50516 43494
rect 50540 43492 50596 43494
rect 53194 45464 53250 45520
rect 50300 42458 50356 42460
rect 50380 42458 50436 42460
rect 50460 42458 50516 42460
rect 50540 42458 50596 42460
rect 50300 42406 50346 42458
rect 50346 42406 50356 42458
rect 50380 42406 50410 42458
rect 50410 42406 50422 42458
rect 50422 42406 50436 42458
rect 50460 42406 50474 42458
rect 50474 42406 50486 42458
rect 50486 42406 50516 42458
rect 50540 42406 50550 42458
rect 50550 42406 50596 42458
rect 50300 42404 50356 42406
rect 50380 42404 50436 42406
rect 50460 42404 50516 42406
rect 50540 42404 50596 42406
rect 50300 41370 50356 41372
rect 50380 41370 50436 41372
rect 50460 41370 50516 41372
rect 50540 41370 50596 41372
rect 50300 41318 50346 41370
rect 50346 41318 50356 41370
rect 50380 41318 50410 41370
rect 50410 41318 50422 41370
rect 50422 41318 50436 41370
rect 50460 41318 50474 41370
rect 50474 41318 50486 41370
rect 50486 41318 50516 41370
rect 50540 41318 50550 41370
rect 50550 41318 50596 41370
rect 50300 41316 50356 41318
rect 50380 41316 50436 41318
rect 50460 41316 50516 41318
rect 50540 41316 50596 41318
rect 50300 40282 50356 40284
rect 50380 40282 50436 40284
rect 50460 40282 50516 40284
rect 50540 40282 50596 40284
rect 50300 40230 50346 40282
rect 50346 40230 50356 40282
rect 50380 40230 50410 40282
rect 50410 40230 50422 40282
rect 50422 40230 50436 40282
rect 50460 40230 50474 40282
rect 50474 40230 50486 40282
rect 50486 40230 50516 40282
rect 50540 40230 50550 40282
rect 50550 40230 50596 40282
rect 50300 40228 50356 40230
rect 50380 40228 50436 40230
rect 50460 40228 50516 40230
rect 50540 40228 50596 40230
rect 50300 39194 50356 39196
rect 50380 39194 50436 39196
rect 50460 39194 50516 39196
rect 50540 39194 50596 39196
rect 50300 39142 50346 39194
rect 50346 39142 50356 39194
rect 50380 39142 50410 39194
rect 50410 39142 50422 39194
rect 50422 39142 50436 39194
rect 50460 39142 50474 39194
rect 50474 39142 50486 39194
rect 50486 39142 50516 39194
rect 50540 39142 50550 39194
rect 50550 39142 50596 39194
rect 50300 39140 50356 39142
rect 50380 39140 50436 39142
rect 50460 39140 50516 39142
rect 50540 39140 50596 39142
rect 50300 38106 50356 38108
rect 50380 38106 50436 38108
rect 50460 38106 50516 38108
rect 50540 38106 50596 38108
rect 50300 38054 50346 38106
rect 50346 38054 50356 38106
rect 50380 38054 50410 38106
rect 50410 38054 50422 38106
rect 50422 38054 50436 38106
rect 50460 38054 50474 38106
rect 50474 38054 50486 38106
rect 50486 38054 50516 38106
rect 50540 38054 50550 38106
rect 50550 38054 50596 38106
rect 50300 38052 50356 38054
rect 50380 38052 50436 38054
rect 50460 38052 50516 38054
rect 50540 38052 50596 38054
rect 50300 37018 50356 37020
rect 50380 37018 50436 37020
rect 50460 37018 50516 37020
rect 50540 37018 50596 37020
rect 50300 36966 50346 37018
rect 50346 36966 50356 37018
rect 50380 36966 50410 37018
rect 50410 36966 50422 37018
rect 50422 36966 50436 37018
rect 50460 36966 50474 37018
rect 50474 36966 50486 37018
rect 50486 36966 50516 37018
rect 50540 36966 50550 37018
rect 50550 36966 50596 37018
rect 50300 36964 50356 36966
rect 50380 36964 50436 36966
rect 50460 36964 50516 36966
rect 50540 36964 50596 36966
rect 50300 35930 50356 35932
rect 50380 35930 50436 35932
rect 50460 35930 50516 35932
rect 50540 35930 50596 35932
rect 50300 35878 50346 35930
rect 50346 35878 50356 35930
rect 50380 35878 50410 35930
rect 50410 35878 50422 35930
rect 50422 35878 50436 35930
rect 50460 35878 50474 35930
rect 50474 35878 50486 35930
rect 50486 35878 50516 35930
rect 50540 35878 50550 35930
rect 50550 35878 50596 35930
rect 50300 35876 50356 35878
rect 50380 35876 50436 35878
rect 50460 35876 50516 35878
rect 50540 35876 50596 35878
rect 50300 34842 50356 34844
rect 50380 34842 50436 34844
rect 50460 34842 50516 34844
rect 50540 34842 50596 34844
rect 50300 34790 50346 34842
rect 50346 34790 50356 34842
rect 50380 34790 50410 34842
rect 50410 34790 50422 34842
rect 50422 34790 50436 34842
rect 50460 34790 50474 34842
rect 50474 34790 50486 34842
rect 50486 34790 50516 34842
rect 50540 34790 50550 34842
rect 50550 34790 50596 34842
rect 50300 34788 50356 34790
rect 50380 34788 50436 34790
rect 50460 34788 50516 34790
rect 50540 34788 50596 34790
rect 50300 33754 50356 33756
rect 50380 33754 50436 33756
rect 50460 33754 50516 33756
rect 50540 33754 50596 33756
rect 50300 33702 50346 33754
rect 50346 33702 50356 33754
rect 50380 33702 50410 33754
rect 50410 33702 50422 33754
rect 50422 33702 50436 33754
rect 50460 33702 50474 33754
rect 50474 33702 50486 33754
rect 50486 33702 50516 33754
rect 50540 33702 50550 33754
rect 50550 33702 50596 33754
rect 50300 33700 50356 33702
rect 50380 33700 50436 33702
rect 50460 33700 50516 33702
rect 50540 33700 50596 33702
rect 50300 32666 50356 32668
rect 50380 32666 50436 32668
rect 50460 32666 50516 32668
rect 50540 32666 50596 32668
rect 50300 32614 50346 32666
rect 50346 32614 50356 32666
rect 50380 32614 50410 32666
rect 50410 32614 50422 32666
rect 50422 32614 50436 32666
rect 50460 32614 50474 32666
rect 50474 32614 50486 32666
rect 50486 32614 50516 32666
rect 50540 32614 50550 32666
rect 50550 32614 50596 32666
rect 50300 32612 50356 32614
rect 50380 32612 50436 32614
rect 50460 32612 50516 32614
rect 50540 32612 50596 32614
rect 50300 31578 50356 31580
rect 50380 31578 50436 31580
rect 50460 31578 50516 31580
rect 50540 31578 50596 31580
rect 50300 31526 50346 31578
rect 50346 31526 50356 31578
rect 50380 31526 50410 31578
rect 50410 31526 50422 31578
rect 50422 31526 50436 31578
rect 50460 31526 50474 31578
rect 50474 31526 50486 31578
rect 50486 31526 50516 31578
rect 50540 31526 50550 31578
rect 50550 31526 50596 31578
rect 50300 31524 50356 31526
rect 50380 31524 50436 31526
rect 50460 31524 50516 31526
rect 50540 31524 50596 31526
rect 50300 30490 50356 30492
rect 50380 30490 50436 30492
rect 50460 30490 50516 30492
rect 50540 30490 50596 30492
rect 50300 30438 50346 30490
rect 50346 30438 50356 30490
rect 50380 30438 50410 30490
rect 50410 30438 50422 30490
rect 50422 30438 50436 30490
rect 50460 30438 50474 30490
rect 50474 30438 50486 30490
rect 50486 30438 50516 30490
rect 50540 30438 50550 30490
rect 50550 30438 50596 30490
rect 50300 30436 50356 30438
rect 50380 30436 50436 30438
rect 50460 30436 50516 30438
rect 50540 30436 50596 30438
rect 50300 29402 50356 29404
rect 50380 29402 50436 29404
rect 50460 29402 50516 29404
rect 50540 29402 50596 29404
rect 50300 29350 50346 29402
rect 50346 29350 50356 29402
rect 50380 29350 50410 29402
rect 50410 29350 50422 29402
rect 50422 29350 50436 29402
rect 50460 29350 50474 29402
rect 50474 29350 50486 29402
rect 50486 29350 50516 29402
rect 50540 29350 50550 29402
rect 50550 29350 50596 29402
rect 50300 29348 50356 29350
rect 50380 29348 50436 29350
rect 50460 29348 50516 29350
rect 50540 29348 50596 29350
rect 50300 28314 50356 28316
rect 50380 28314 50436 28316
rect 50460 28314 50516 28316
rect 50540 28314 50596 28316
rect 50300 28262 50346 28314
rect 50346 28262 50356 28314
rect 50380 28262 50410 28314
rect 50410 28262 50422 28314
rect 50422 28262 50436 28314
rect 50460 28262 50474 28314
rect 50474 28262 50486 28314
rect 50486 28262 50516 28314
rect 50540 28262 50550 28314
rect 50550 28262 50596 28314
rect 50300 28260 50356 28262
rect 50380 28260 50436 28262
rect 50460 28260 50516 28262
rect 50540 28260 50596 28262
rect 50300 27226 50356 27228
rect 50380 27226 50436 27228
rect 50460 27226 50516 27228
rect 50540 27226 50596 27228
rect 50300 27174 50346 27226
rect 50346 27174 50356 27226
rect 50380 27174 50410 27226
rect 50410 27174 50422 27226
rect 50422 27174 50436 27226
rect 50460 27174 50474 27226
rect 50474 27174 50486 27226
rect 50486 27174 50516 27226
rect 50540 27174 50550 27226
rect 50550 27174 50596 27226
rect 50300 27172 50356 27174
rect 50380 27172 50436 27174
rect 50460 27172 50516 27174
rect 50540 27172 50596 27174
rect 50300 26138 50356 26140
rect 50380 26138 50436 26140
rect 50460 26138 50516 26140
rect 50540 26138 50596 26140
rect 50300 26086 50346 26138
rect 50346 26086 50356 26138
rect 50380 26086 50410 26138
rect 50410 26086 50422 26138
rect 50422 26086 50436 26138
rect 50460 26086 50474 26138
rect 50474 26086 50486 26138
rect 50486 26086 50516 26138
rect 50540 26086 50550 26138
rect 50550 26086 50596 26138
rect 50300 26084 50356 26086
rect 50380 26084 50436 26086
rect 50460 26084 50516 26086
rect 50540 26084 50596 26086
rect 50300 25050 50356 25052
rect 50380 25050 50436 25052
rect 50460 25050 50516 25052
rect 50540 25050 50596 25052
rect 50300 24998 50346 25050
rect 50346 24998 50356 25050
rect 50380 24998 50410 25050
rect 50410 24998 50422 25050
rect 50422 24998 50436 25050
rect 50460 24998 50474 25050
rect 50474 24998 50486 25050
rect 50486 24998 50516 25050
rect 50540 24998 50550 25050
rect 50550 24998 50596 25050
rect 50300 24996 50356 24998
rect 50380 24996 50436 24998
rect 50460 24996 50516 24998
rect 50540 24996 50596 24998
rect 50300 23962 50356 23964
rect 50380 23962 50436 23964
rect 50460 23962 50516 23964
rect 50540 23962 50596 23964
rect 50300 23910 50346 23962
rect 50346 23910 50356 23962
rect 50380 23910 50410 23962
rect 50410 23910 50422 23962
rect 50422 23910 50436 23962
rect 50460 23910 50474 23962
rect 50474 23910 50486 23962
rect 50486 23910 50516 23962
rect 50540 23910 50550 23962
rect 50550 23910 50596 23962
rect 50300 23908 50356 23910
rect 50380 23908 50436 23910
rect 50460 23908 50516 23910
rect 50540 23908 50596 23910
rect 58162 46996 58164 47016
rect 58164 46996 58216 47016
rect 58216 46996 58218 47016
rect 58162 46960 58218 46996
rect 58162 42200 58218 42256
rect 58162 32000 58218 32056
rect 57702 29280 57758 29336
rect 50300 22874 50356 22876
rect 50380 22874 50436 22876
rect 50460 22874 50516 22876
rect 50540 22874 50596 22876
rect 50300 22822 50346 22874
rect 50346 22822 50356 22874
rect 50380 22822 50410 22874
rect 50410 22822 50422 22874
rect 50422 22822 50436 22874
rect 50460 22822 50474 22874
rect 50474 22822 50486 22874
rect 50486 22822 50516 22874
rect 50540 22822 50550 22874
rect 50550 22822 50596 22874
rect 50300 22820 50356 22822
rect 50380 22820 50436 22822
rect 50460 22820 50516 22822
rect 50540 22820 50596 22822
rect 50300 21786 50356 21788
rect 50380 21786 50436 21788
rect 50460 21786 50516 21788
rect 50540 21786 50596 21788
rect 50300 21734 50346 21786
rect 50346 21734 50356 21786
rect 50380 21734 50410 21786
rect 50410 21734 50422 21786
rect 50422 21734 50436 21786
rect 50460 21734 50474 21786
rect 50474 21734 50486 21786
rect 50486 21734 50516 21786
rect 50540 21734 50550 21786
rect 50550 21734 50596 21786
rect 50300 21732 50356 21734
rect 50380 21732 50436 21734
rect 50460 21732 50516 21734
rect 50540 21732 50596 21734
rect 50300 20698 50356 20700
rect 50380 20698 50436 20700
rect 50460 20698 50516 20700
rect 50540 20698 50596 20700
rect 50300 20646 50346 20698
rect 50346 20646 50356 20698
rect 50380 20646 50410 20698
rect 50410 20646 50422 20698
rect 50422 20646 50436 20698
rect 50460 20646 50474 20698
rect 50474 20646 50486 20698
rect 50486 20646 50516 20698
rect 50540 20646 50550 20698
rect 50550 20646 50596 20698
rect 50300 20644 50356 20646
rect 50380 20644 50436 20646
rect 50460 20644 50516 20646
rect 50540 20644 50596 20646
rect 50300 19610 50356 19612
rect 50380 19610 50436 19612
rect 50460 19610 50516 19612
rect 50540 19610 50596 19612
rect 50300 19558 50346 19610
rect 50346 19558 50356 19610
rect 50380 19558 50410 19610
rect 50410 19558 50422 19610
rect 50422 19558 50436 19610
rect 50460 19558 50474 19610
rect 50474 19558 50486 19610
rect 50486 19558 50516 19610
rect 50540 19558 50550 19610
rect 50550 19558 50596 19610
rect 50300 19556 50356 19558
rect 50380 19556 50436 19558
rect 50460 19556 50516 19558
rect 50540 19556 50596 19558
rect 50300 18522 50356 18524
rect 50380 18522 50436 18524
rect 50460 18522 50516 18524
rect 50540 18522 50596 18524
rect 50300 18470 50346 18522
rect 50346 18470 50356 18522
rect 50380 18470 50410 18522
rect 50410 18470 50422 18522
rect 50422 18470 50436 18522
rect 50460 18470 50474 18522
rect 50474 18470 50486 18522
rect 50486 18470 50516 18522
rect 50540 18470 50550 18522
rect 50550 18470 50596 18522
rect 50300 18468 50356 18470
rect 50380 18468 50436 18470
rect 50460 18468 50516 18470
rect 50540 18468 50596 18470
rect 50300 17434 50356 17436
rect 50380 17434 50436 17436
rect 50460 17434 50516 17436
rect 50540 17434 50596 17436
rect 50300 17382 50346 17434
rect 50346 17382 50356 17434
rect 50380 17382 50410 17434
rect 50410 17382 50422 17434
rect 50422 17382 50436 17434
rect 50460 17382 50474 17434
rect 50474 17382 50486 17434
rect 50486 17382 50516 17434
rect 50540 17382 50550 17434
rect 50550 17382 50596 17434
rect 50300 17380 50356 17382
rect 50380 17380 50436 17382
rect 50460 17380 50516 17382
rect 50540 17380 50596 17382
rect 50300 16346 50356 16348
rect 50380 16346 50436 16348
rect 50460 16346 50516 16348
rect 50540 16346 50596 16348
rect 50300 16294 50346 16346
rect 50346 16294 50356 16346
rect 50380 16294 50410 16346
rect 50410 16294 50422 16346
rect 50422 16294 50436 16346
rect 50460 16294 50474 16346
rect 50474 16294 50486 16346
rect 50486 16294 50516 16346
rect 50540 16294 50550 16346
rect 50550 16294 50596 16346
rect 50300 16292 50356 16294
rect 50380 16292 50436 16294
rect 50460 16292 50516 16294
rect 50540 16292 50596 16294
rect 50300 15258 50356 15260
rect 50380 15258 50436 15260
rect 50460 15258 50516 15260
rect 50540 15258 50596 15260
rect 50300 15206 50346 15258
rect 50346 15206 50356 15258
rect 50380 15206 50410 15258
rect 50410 15206 50422 15258
rect 50422 15206 50436 15258
rect 50460 15206 50474 15258
rect 50474 15206 50486 15258
rect 50486 15206 50516 15258
rect 50540 15206 50550 15258
rect 50550 15206 50596 15258
rect 50300 15204 50356 15206
rect 50380 15204 50436 15206
rect 50460 15204 50516 15206
rect 50540 15204 50596 15206
rect 50300 14170 50356 14172
rect 50380 14170 50436 14172
rect 50460 14170 50516 14172
rect 50540 14170 50596 14172
rect 50300 14118 50346 14170
rect 50346 14118 50356 14170
rect 50380 14118 50410 14170
rect 50410 14118 50422 14170
rect 50422 14118 50436 14170
rect 50460 14118 50474 14170
rect 50474 14118 50486 14170
rect 50486 14118 50516 14170
rect 50540 14118 50550 14170
rect 50550 14118 50596 14170
rect 50300 14116 50356 14118
rect 50380 14116 50436 14118
rect 50460 14116 50516 14118
rect 50540 14116 50596 14118
rect 50300 13082 50356 13084
rect 50380 13082 50436 13084
rect 50460 13082 50516 13084
rect 50540 13082 50596 13084
rect 50300 13030 50346 13082
rect 50346 13030 50356 13082
rect 50380 13030 50410 13082
rect 50410 13030 50422 13082
rect 50422 13030 50436 13082
rect 50460 13030 50474 13082
rect 50474 13030 50486 13082
rect 50486 13030 50516 13082
rect 50540 13030 50550 13082
rect 50550 13030 50596 13082
rect 50300 13028 50356 13030
rect 50380 13028 50436 13030
rect 50460 13028 50516 13030
rect 50540 13028 50596 13030
rect 50300 11994 50356 11996
rect 50380 11994 50436 11996
rect 50460 11994 50516 11996
rect 50540 11994 50596 11996
rect 50300 11942 50346 11994
rect 50346 11942 50356 11994
rect 50380 11942 50410 11994
rect 50410 11942 50422 11994
rect 50422 11942 50436 11994
rect 50460 11942 50474 11994
rect 50474 11942 50486 11994
rect 50486 11942 50516 11994
rect 50540 11942 50550 11994
rect 50550 11942 50596 11994
rect 50300 11940 50356 11942
rect 50380 11940 50436 11942
rect 50460 11940 50516 11942
rect 50540 11940 50596 11942
rect 50300 10906 50356 10908
rect 50380 10906 50436 10908
rect 50460 10906 50516 10908
rect 50540 10906 50596 10908
rect 50300 10854 50346 10906
rect 50346 10854 50356 10906
rect 50380 10854 50410 10906
rect 50410 10854 50422 10906
rect 50422 10854 50436 10906
rect 50460 10854 50474 10906
rect 50474 10854 50486 10906
rect 50486 10854 50516 10906
rect 50540 10854 50550 10906
rect 50550 10854 50596 10906
rect 50300 10852 50356 10854
rect 50380 10852 50436 10854
rect 50460 10852 50516 10854
rect 50540 10852 50596 10854
rect 50300 9818 50356 9820
rect 50380 9818 50436 9820
rect 50460 9818 50516 9820
rect 50540 9818 50596 9820
rect 50300 9766 50346 9818
rect 50346 9766 50356 9818
rect 50380 9766 50410 9818
rect 50410 9766 50422 9818
rect 50422 9766 50436 9818
rect 50460 9766 50474 9818
rect 50474 9766 50486 9818
rect 50486 9766 50516 9818
rect 50540 9766 50550 9818
rect 50550 9766 50596 9818
rect 50300 9764 50356 9766
rect 50380 9764 50436 9766
rect 50460 9764 50516 9766
rect 50540 9764 50596 9766
rect 50300 8730 50356 8732
rect 50380 8730 50436 8732
rect 50460 8730 50516 8732
rect 50540 8730 50596 8732
rect 50300 8678 50346 8730
rect 50346 8678 50356 8730
rect 50380 8678 50410 8730
rect 50410 8678 50422 8730
rect 50422 8678 50436 8730
rect 50460 8678 50474 8730
rect 50474 8678 50486 8730
rect 50486 8678 50516 8730
rect 50540 8678 50550 8730
rect 50550 8678 50596 8730
rect 50300 8676 50356 8678
rect 50380 8676 50436 8678
rect 50460 8676 50516 8678
rect 50540 8676 50596 8678
rect 50300 7642 50356 7644
rect 50380 7642 50436 7644
rect 50460 7642 50516 7644
rect 50540 7642 50596 7644
rect 50300 7590 50346 7642
rect 50346 7590 50356 7642
rect 50380 7590 50410 7642
rect 50410 7590 50422 7642
rect 50422 7590 50436 7642
rect 50460 7590 50474 7642
rect 50474 7590 50486 7642
rect 50486 7590 50516 7642
rect 50540 7590 50550 7642
rect 50550 7590 50596 7642
rect 50300 7588 50356 7590
rect 50380 7588 50436 7590
rect 50460 7588 50516 7590
rect 50540 7588 50596 7590
rect 50300 6554 50356 6556
rect 50380 6554 50436 6556
rect 50460 6554 50516 6556
rect 50540 6554 50596 6556
rect 50300 6502 50346 6554
rect 50346 6502 50356 6554
rect 50380 6502 50410 6554
rect 50410 6502 50422 6554
rect 50422 6502 50436 6554
rect 50460 6502 50474 6554
rect 50474 6502 50486 6554
rect 50486 6502 50516 6554
rect 50540 6502 50550 6554
rect 50550 6502 50596 6554
rect 50300 6500 50356 6502
rect 50380 6500 50436 6502
rect 50460 6500 50516 6502
rect 50540 6500 50596 6502
rect 50300 5466 50356 5468
rect 50380 5466 50436 5468
rect 50460 5466 50516 5468
rect 50540 5466 50596 5468
rect 50300 5414 50346 5466
rect 50346 5414 50356 5466
rect 50380 5414 50410 5466
rect 50410 5414 50422 5466
rect 50422 5414 50436 5466
rect 50460 5414 50474 5466
rect 50474 5414 50486 5466
rect 50486 5414 50516 5466
rect 50540 5414 50550 5466
rect 50550 5414 50596 5466
rect 50300 5412 50356 5414
rect 50380 5412 50436 5414
rect 50460 5412 50516 5414
rect 50540 5412 50596 5414
rect 50300 4378 50356 4380
rect 50380 4378 50436 4380
rect 50460 4378 50516 4380
rect 50540 4378 50596 4380
rect 50300 4326 50346 4378
rect 50346 4326 50356 4378
rect 50380 4326 50410 4378
rect 50410 4326 50422 4378
rect 50422 4326 50436 4378
rect 50460 4326 50474 4378
rect 50474 4326 50486 4378
rect 50486 4326 50516 4378
rect 50540 4326 50550 4378
rect 50550 4326 50596 4378
rect 50300 4324 50356 4326
rect 50380 4324 50436 4326
rect 50460 4324 50516 4326
rect 50540 4324 50596 4326
rect 50300 3290 50356 3292
rect 50380 3290 50436 3292
rect 50460 3290 50516 3292
rect 50540 3290 50596 3292
rect 50300 3238 50346 3290
rect 50346 3238 50356 3290
rect 50380 3238 50410 3290
rect 50410 3238 50422 3290
rect 50422 3238 50436 3290
rect 50460 3238 50474 3290
rect 50474 3238 50486 3290
rect 50486 3238 50516 3290
rect 50540 3238 50550 3290
rect 50550 3238 50596 3290
rect 50300 3236 50356 3238
rect 50380 3236 50436 3238
rect 50460 3236 50516 3238
rect 50540 3236 50596 3238
rect 50300 2202 50356 2204
rect 50380 2202 50436 2204
rect 50460 2202 50516 2204
rect 50540 2202 50596 2204
rect 50300 2150 50346 2202
rect 50346 2150 50356 2202
rect 50380 2150 50410 2202
rect 50410 2150 50422 2202
rect 50422 2150 50436 2202
rect 50460 2150 50474 2202
rect 50474 2150 50486 2202
rect 50486 2150 50516 2202
rect 50540 2150 50550 2202
rect 50550 2150 50596 2202
rect 50300 2148 50356 2150
rect 50380 2148 50436 2150
rect 50460 2148 50516 2150
rect 50540 2148 50596 2150
rect 58162 24520 58218 24576
rect 58162 19080 58218 19136
rect 58162 11600 58218 11656
rect 58162 8900 58218 8936
rect 58162 8880 58164 8900
rect 58164 8880 58216 8900
rect 58216 8880 58218 8900
rect 57886 1400 57942 1456
<< metal3 >>
rect 0 57748 800 57988
rect 19568 57696 19888 57697
rect 19568 57632 19576 57696
rect 19640 57632 19656 57696
rect 19720 57632 19736 57696
rect 19800 57632 19816 57696
rect 19880 57632 19888 57696
rect 19568 57631 19888 57632
rect 50288 57696 50608 57697
rect 50288 57632 50296 57696
rect 50360 57632 50376 57696
rect 50440 57632 50456 57696
rect 50520 57632 50536 57696
rect 50600 57632 50608 57696
rect 50288 57631 50608 57632
rect 4208 57152 4528 57153
rect 4208 57088 4216 57152
rect 4280 57088 4296 57152
rect 4360 57088 4376 57152
rect 4440 57088 4456 57152
rect 4520 57088 4528 57152
rect 4208 57087 4528 57088
rect 34928 57152 35248 57153
rect 34928 57088 34936 57152
rect 35000 57088 35016 57152
rect 35080 57088 35096 57152
rect 35160 57088 35176 57152
rect 35240 57088 35248 57152
rect 34928 57087 35248 57088
rect 59200 57068 60000 57308
rect 19568 56608 19888 56609
rect 19568 56544 19576 56608
rect 19640 56544 19656 56608
rect 19720 56544 19736 56608
rect 19800 56544 19816 56608
rect 19880 56544 19888 56608
rect 19568 56543 19888 56544
rect 50288 56608 50608 56609
rect 50288 56544 50296 56608
rect 50360 56544 50376 56608
rect 50440 56544 50456 56608
rect 50520 56544 50536 56608
rect 50600 56544 50608 56608
rect 50288 56543 50608 56544
rect 4208 56064 4528 56065
rect 4208 56000 4216 56064
rect 4280 56000 4296 56064
rect 4360 56000 4376 56064
rect 4440 56000 4456 56064
rect 4520 56000 4528 56064
rect 4208 55999 4528 56000
rect 34928 56064 35248 56065
rect 34928 56000 34936 56064
rect 35000 56000 35016 56064
rect 35080 56000 35096 56064
rect 35160 56000 35176 56064
rect 35240 56000 35248 56064
rect 34928 55999 35248 56000
rect 19568 55520 19888 55521
rect 19568 55456 19576 55520
rect 19640 55456 19656 55520
rect 19720 55456 19736 55520
rect 19800 55456 19816 55520
rect 19880 55456 19888 55520
rect 19568 55455 19888 55456
rect 50288 55520 50608 55521
rect 50288 55456 50296 55520
rect 50360 55456 50376 55520
rect 50440 55456 50456 55520
rect 50520 55456 50536 55520
rect 50600 55456 50608 55520
rect 50288 55455 50608 55456
rect 0 55178 800 55268
rect 2773 55178 2839 55181
rect 0 55176 2839 55178
rect 0 55120 2778 55176
rect 2834 55120 2839 55176
rect 0 55118 2839 55120
rect 0 55028 800 55118
rect 2773 55115 2839 55118
rect 4208 54976 4528 54977
rect 4208 54912 4216 54976
rect 4280 54912 4296 54976
rect 4360 54912 4376 54976
rect 4440 54912 4456 54976
rect 4520 54912 4528 54976
rect 4208 54911 4528 54912
rect 34928 54976 35248 54977
rect 34928 54912 34936 54976
rect 35000 54912 35016 54976
rect 35080 54912 35096 54976
rect 35160 54912 35176 54976
rect 35240 54912 35248 54976
rect 34928 54911 35248 54912
rect 19568 54432 19888 54433
rect 19568 54368 19576 54432
rect 19640 54368 19656 54432
rect 19720 54368 19736 54432
rect 19800 54368 19816 54432
rect 19880 54368 19888 54432
rect 19568 54367 19888 54368
rect 50288 54432 50608 54433
rect 50288 54368 50296 54432
rect 50360 54368 50376 54432
rect 50440 54368 50456 54432
rect 50520 54368 50536 54432
rect 50600 54368 50608 54432
rect 50288 54367 50608 54368
rect 59200 54348 60000 54588
rect 4208 53888 4528 53889
rect 4208 53824 4216 53888
rect 4280 53824 4296 53888
rect 4360 53824 4376 53888
rect 4440 53824 4456 53888
rect 4520 53824 4528 53888
rect 4208 53823 4528 53824
rect 34928 53888 35248 53889
rect 34928 53824 34936 53888
rect 35000 53824 35016 53888
rect 35080 53824 35096 53888
rect 35160 53824 35176 53888
rect 35240 53824 35248 53888
rect 34928 53823 35248 53824
rect 19568 53344 19888 53345
rect 19568 53280 19576 53344
rect 19640 53280 19656 53344
rect 19720 53280 19736 53344
rect 19800 53280 19816 53344
rect 19880 53280 19888 53344
rect 19568 53279 19888 53280
rect 50288 53344 50608 53345
rect 50288 53280 50296 53344
rect 50360 53280 50376 53344
rect 50440 53280 50456 53344
rect 50520 53280 50536 53344
rect 50600 53280 50608 53344
rect 50288 53279 50608 53280
rect 4208 52800 4528 52801
rect 4208 52736 4216 52800
rect 4280 52736 4296 52800
rect 4360 52736 4376 52800
rect 4440 52736 4456 52800
rect 4520 52736 4528 52800
rect 4208 52735 4528 52736
rect 34928 52800 35248 52801
rect 34928 52736 34936 52800
rect 35000 52736 35016 52800
rect 35080 52736 35096 52800
rect 35160 52736 35176 52800
rect 35240 52736 35248 52800
rect 34928 52735 35248 52736
rect 0 52308 800 52548
rect 19568 52256 19888 52257
rect 19568 52192 19576 52256
rect 19640 52192 19656 52256
rect 19720 52192 19736 52256
rect 19800 52192 19816 52256
rect 19880 52192 19888 52256
rect 19568 52191 19888 52192
rect 50288 52256 50608 52257
rect 50288 52192 50296 52256
rect 50360 52192 50376 52256
rect 50440 52192 50456 52256
rect 50520 52192 50536 52256
rect 50600 52192 50608 52256
rect 50288 52191 50608 52192
rect 4208 51712 4528 51713
rect 4208 51648 4216 51712
rect 4280 51648 4296 51712
rect 4360 51648 4376 51712
rect 4440 51648 4456 51712
rect 4520 51648 4528 51712
rect 4208 51647 4528 51648
rect 34928 51712 35248 51713
rect 34928 51648 34936 51712
rect 35000 51648 35016 51712
rect 35080 51648 35096 51712
rect 35160 51648 35176 51712
rect 35240 51648 35248 51712
rect 34928 51647 35248 51648
rect 59200 51628 60000 51868
rect 19568 51168 19888 51169
rect 19568 51104 19576 51168
rect 19640 51104 19656 51168
rect 19720 51104 19736 51168
rect 19800 51104 19816 51168
rect 19880 51104 19888 51168
rect 19568 51103 19888 51104
rect 50288 51168 50608 51169
rect 50288 51104 50296 51168
rect 50360 51104 50376 51168
rect 50440 51104 50456 51168
rect 50520 51104 50536 51168
rect 50600 51104 50608 51168
rect 50288 51103 50608 51104
rect 4208 50624 4528 50625
rect 4208 50560 4216 50624
rect 4280 50560 4296 50624
rect 4360 50560 4376 50624
rect 4440 50560 4456 50624
rect 4520 50560 4528 50624
rect 4208 50559 4528 50560
rect 34928 50624 35248 50625
rect 34928 50560 34936 50624
rect 35000 50560 35016 50624
rect 35080 50560 35096 50624
rect 35160 50560 35176 50624
rect 35240 50560 35248 50624
rect 34928 50559 35248 50560
rect 0 50418 800 50508
rect 2773 50418 2839 50421
rect 0 50416 2839 50418
rect 0 50360 2778 50416
rect 2834 50360 2839 50416
rect 0 50358 2839 50360
rect 0 50268 800 50358
rect 2773 50355 2839 50358
rect 19568 50080 19888 50081
rect 19568 50016 19576 50080
rect 19640 50016 19656 50080
rect 19720 50016 19736 50080
rect 19800 50016 19816 50080
rect 19880 50016 19888 50080
rect 19568 50015 19888 50016
rect 50288 50080 50608 50081
rect 50288 50016 50296 50080
rect 50360 50016 50376 50080
rect 50440 50016 50456 50080
rect 50520 50016 50536 50080
rect 50600 50016 50608 50080
rect 50288 50015 50608 50016
rect 59200 49588 60000 49828
rect 4208 49536 4528 49537
rect 4208 49472 4216 49536
rect 4280 49472 4296 49536
rect 4360 49472 4376 49536
rect 4440 49472 4456 49536
rect 4520 49472 4528 49536
rect 4208 49471 4528 49472
rect 34928 49536 35248 49537
rect 34928 49472 34936 49536
rect 35000 49472 35016 49536
rect 35080 49472 35096 49536
rect 35160 49472 35176 49536
rect 35240 49472 35248 49536
rect 34928 49471 35248 49472
rect 19568 48992 19888 48993
rect 19568 48928 19576 48992
rect 19640 48928 19656 48992
rect 19720 48928 19736 48992
rect 19800 48928 19816 48992
rect 19880 48928 19888 48992
rect 19568 48927 19888 48928
rect 50288 48992 50608 48993
rect 50288 48928 50296 48992
rect 50360 48928 50376 48992
rect 50440 48928 50456 48992
rect 50520 48928 50536 48992
rect 50600 48928 50608 48992
rect 50288 48927 50608 48928
rect 4208 48448 4528 48449
rect 4208 48384 4216 48448
rect 4280 48384 4296 48448
rect 4360 48384 4376 48448
rect 4440 48384 4456 48448
rect 4520 48384 4528 48448
rect 4208 48383 4528 48384
rect 34928 48448 35248 48449
rect 34928 48384 34936 48448
rect 35000 48384 35016 48448
rect 35080 48384 35096 48448
rect 35160 48384 35176 48448
rect 35240 48384 35248 48448
rect 34928 48383 35248 48384
rect 19568 47904 19888 47905
rect 19568 47840 19576 47904
rect 19640 47840 19656 47904
rect 19720 47840 19736 47904
rect 19800 47840 19816 47904
rect 19880 47840 19888 47904
rect 19568 47839 19888 47840
rect 50288 47904 50608 47905
rect 50288 47840 50296 47904
rect 50360 47840 50376 47904
rect 50440 47840 50456 47904
rect 50520 47840 50536 47904
rect 50600 47840 50608 47904
rect 50288 47839 50608 47840
rect 0 47698 800 47788
rect 2773 47698 2839 47701
rect 0 47696 2839 47698
rect 0 47640 2778 47696
rect 2834 47640 2839 47696
rect 0 47638 2839 47640
rect 0 47548 800 47638
rect 2773 47635 2839 47638
rect 4208 47360 4528 47361
rect 4208 47296 4216 47360
rect 4280 47296 4296 47360
rect 4360 47296 4376 47360
rect 4440 47296 4456 47360
rect 4520 47296 4528 47360
rect 4208 47295 4528 47296
rect 34928 47360 35248 47361
rect 34928 47296 34936 47360
rect 35000 47296 35016 47360
rect 35080 47296 35096 47360
rect 35160 47296 35176 47360
rect 35240 47296 35248 47360
rect 34928 47295 35248 47296
rect 58157 47018 58223 47021
rect 59200 47018 60000 47108
rect 58157 47016 60000 47018
rect 58157 46960 58162 47016
rect 58218 46960 60000 47016
rect 58157 46958 60000 46960
rect 58157 46955 58223 46958
rect 59200 46868 60000 46958
rect 19568 46816 19888 46817
rect 19568 46752 19576 46816
rect 19640 46752 19656 46816
rect 19720 46752 19736 46816
rect 19800 46752 19816 46816
rect 19880 46752 19888 46816
rect 19568 46751 19888 46752
rect 50288 46816 50608 46817
rect 50288 46752 50296 46816
rect 50360 46752 50376 46816
rect 50440 46752 50456 46816
rect 50520 46752 50536 46816
rect 50600 46752 50608 46816
rect 50288 46751 50608 46752
rect 4208 46272 4528 46273
rect 4208 46208 4216 46272
rect 4280 46208 4296 46272
rect 4360 46208 4376 46272
rect 4440 46208 4456 46272
rect 4520 46208 4528 46272
rect 4208 46207 4528 46208
rect 34928 46272 35248 46273
rect 34928 46208 34936 46272
rect 35000 46208 35016 46272
rect 35080 46208 35096 46272
rect 35160 46208 35176 46272
rect 35240 46208 35248 46272
rect 34928 46207 35248 46208
rect 19568 45728 19888 45729
rect 19568 45664 19576 45728
rect 19640 45664 19656 45728
rect 19720 45664 19736 45728
rect 19800 45664 19816 45728
rect 19880 45664 19888 45728
rect 19568 45663 19888 45664
rect 50288 45728 50608 45729
rect 50288 45664 50296 45728
rect 50360 45664 50376 45728
rect 50440 45664 50456 45728
rect 50520 45664 50536 45728
rect 50600 45664 50608 45728
rect 50288 45663 50608 45664
rect 50981 45522 51047 45525
rect 52637 45522 52703 45525
rect 53189 45522 53255 45525
rect 50981 45520 53255 45522
rect 50981 45464 50986 45520
rect 51042 45464 52642 45520
rect 52698 45464 53194 45520
rect 53250 45464 53255 45520
rect 50981 45462 53255 45464
rect 50981 45459 51047 45462
rect 52637 45459 52703 45462
rect 53189 45459 53255 45462
rect 4208 45184 4528 45185
rect 4208 45120 4216 45184
rect 4280 45120 4296 45184
rect 4360 45120 4376 45184
rect 4440 45120 4456 45184
rect 4520 45120 4528 45184
rect 4208 45119 4528 45120
rect 34928 45184 35248 45185
rect 34928 45120 34936 45184
rect 35000 45120 35016 45184
rect 35080 45120 35096 45184
rect 35160 45120 35176 45184
rect 35240 45120 35248 45184
rect 34928 45119 35248 45120
rect 0 44978 800 45068
rect 2773 44978 2839 44981
rect 0 44976 2839 44978
rect 0 44920 2778 44976
rect 2834 44920 2839 44976
rect 0 44918 2839 44920
rect 0 44828 800 44918
rect 2773 44915 2839 44918
rect 19568 44640 19888 44641
rect 19568 44576 19576 44640
rect 19640 44576 19656 44640
rect 19720 44576 19736 44640
rect 19800 44576 19816 44640
rect 19880 44576 19888 44640
rect 19568 44575 19888 44576
rect 50288 44640 50608 44641
rect 50288 44576 50296 44640
rect 50360 44576 50376 44640
rect 50440 44576 50456 44640
rect 50520 44576 50536 44640
rect 50600 44576 50608 44640
rect 50288 44575 50608 44576
rect 59200 44148 60000 44388
rect 4208 44096 4528 44097
rect 4208 44032 4216 44096
rect 4280 44032 4296 44096
rect 4360 44032 4376 44096
rect 4440 44032 4456 44096
rect 4520 44032 4528 44096
rect 4208 44031 4528 44032
rect 34928 44096 35248 44097
rect 34928 44032 34936 44096
rect 35000 44032 35016 44096
rect 35080 44032 35096 44096
rect 35160 44032 35176 44096
rect 35240 44032 35248 44096
rect 34928 44031 35248 44032
rect 19568 43552 19888 43553
rect 19568 43488 19576 43552
rect 19640 43488 19656 43552
rect 19720 43488 19736 43552
rect 19800 43488 19816 43552
rect 19880 43488 19888 43552
rect 19568 43487 19888 43488
rect 50288 43552 50608 43553
rect 50288 43488 50296 43552
rect 50360 43488 50376 43552
rect 50440 43488 50456 43552
rect 50520 43488 50536 43552
rect 50600 43488 50608 43552
rect 50288 43487 50608 43488
rect 0 42938 800 43028
rect 4208 43008 4528 43009
rect 4208 42944 4216 43008
rect 4280 42944 4296 43008
rect 4360 42944 4376 43008
rect 4440 42944 4456 43008
rect 4520 42944 4528 43008
rect 4208 42943 4528 42944
rect 34928 43008 35248 43009
rect 34928 42944 34936 43008
rect 35000 42944 35016 43008
rect 35080 42944 35096 43008
rect 35160 42944 35176 43008
rect 35240 42944 35248 43008
rect 34928 42943 35248 42944
rect 2773 42938 2839 42941
rect 0 42936 2839 42938
rect 0 42880 2778 42936
rect 2834 42880 2839 42936
rect 0 42878 2839 42880
rect 0 42788 800 42878
rect 2773 42875 2839 42878
rect 19568 42464 19888 42465
rect 19568 42400 19576 42464
rect 19640 42400 19656 42464
rect 19720 42400 19736 42464
rect 19800 42400 19816 42464
rect 19880 42400 19888 42464
rect 19568 42399 19888 42400
rect 50288 42464 50608 42465
rect 50288 42400 50296 42464
rect 50360 42400 50376 42464
rect 50440 42400 50456 42464
rect 50520 42400 50536 42464
rect 50600 42400 50608 42464
rect 50288 42399 50608 42400
rect 58157 42258 58223 42261
rect 59200 42258 60000 42348
rect 58157 42256 60000 42258
rect 58157 42200 58162 42256
rect 58218 42200 60000 42256
rect 58157 42198 60000 42200
rect 58157 42195 58223 42198
rect 59200 42108 60000 42198
rect 4208 41920 4528 41921
rect 4208 41856 4216 41920
rect 4280 41856 4296 41920
rect 4360 41856 4376 41920
rect 4440 41856 4456 41920
rect 4520 41856 4528 41920
rect 4208 41855 4528 41856
rect 34928 41920 35248 41921
rect 34928 41856 34936 41920
rect 35000 41856 35016 41920
rect 35080 41856 35096 41920
rect 35160 41856 35176 41920
rect 35240 41856 35248 41920
rect 34928 41855 35248 41856
rect 19568 41376 19888 41377
rect 19568 41312 19576 41376
rect 19640 41312 19656 41376
rect 19720 41312 19736 41376
rect 19800 41312 19816 41376
rect 19880 41312 19888 41376
rect 19568 41311 19888 41312
rect 50288 41376 50608 41377
rect 50288 41312 50296 41376
rect 50360 41312 50376 41376
rect 50440 41312 50456 41376
rect 50520 41312 50536 41376
rect 50600 41312 50608 41376
rect 50288 41311 50608 41312
rect 4208 40832 4528 40833
rect 4208 40768 4216 40832
rect 4280 40768 4296 40832
rect 4360 40768 4376 40832
rect 4440 40768 4456 40832
rect 4520 40768 4528 40832
rect 4208 40767 4528 40768
rect 34928 40832 35248 40833
rect 34928 40768 34936 40832
rect 35000 40768 35016 40832
rect 35080 40768 35096 40832
rect 35160 40768 35176 40832
rect 35240 40768 35248 40832
rect 34928 40767 35248 40768
rect 0 40068 800 40308
rect 19568 40288 19888 40289
rect 19568 40224 19576 40288
rect 19640 40224 19656 40288
rect 19720 40224 19736 40288
rect 19800 40224 19816 40288
rect 19880 40224 19888 40288
rect 19568 40223 19888 40224
rect 50288 40288 50608 40289
rect 50288 40224 50296 40288
rect 50360 40224 50376 40288
rect 50440 40224 50456 40288
rect 50520 40224 50536 40288
rect 50600 40224 50608 40288
rect 50288 40223 50608 40224
rect 4208 39744 4528 39745
rect 4208 39680 4216 39744
rect 4280 39680 4296 39744
rect 4360 39680 4376 39744
rect 4440 39680 4456 39744
rect 4520 39680 4528 39744
rect 4208 39679 4528 39680
rect 34928 39744 35248 39745
rect 34928 39680 34936 39744
rect 35000 39680 35016 39744
rect 35080 39680 35096 39744
rect 35160 39680 35176 39744
rect 35240 39680 35248 39744
rect 34928 39679 35248 39680
rect 59200 39388 60000 39628
rect 19568 39200 19888 39201
rect 19568 39136 19576 39200
rect 19640 39136 19656 39200
rect 19720 39136 19736 39200
rect 19800 39136 19816 39200
rect 19880 39136 19888 39200
rect 19568 39135 19888 39136
rect 50288 39200 50608 39201
rect 50288 39136 50296 39200
rect 50360 39136 50376 39200
rect 50440 39136 50456 39200
rect 50520 39136 50536 39200
rect 50600 39136 50608 39200
rect 50288 39135 50608 39136
rect 4208 38656 4528 38657
rect 4208 38592 4216 38656
rect 4280 38592 4296 38656
rect 4360 38592 4376 38656
rect 4440 38592 4456 38656
rect 4520 38592 4528 38656
rect 4208 38591 4528 38592
rect 34928 38656 35248 38657
rect 34928 38592 34936 38656
rect 35000 38592 35016 38656
rect 35080 38592 35096 38656
rect 35160 38592 35176 38656
rect 35240 38592 35248 38656
rect 34928 38591 35248 38592
rect 19568 38112 19888 38113
rect 19568 38048 19576 38112
rect 19640 38048 19656 38112
rect 19720 38048 19736 38112
rect 19800 38048 19816 38112
rect 19880 38048 19888 38112
rect 19568 38047 19888 38048
rect 50288 38112 50608 38113
rect 50288 38048 50296 38112
rect 50360 38048 50376 38112
rect 50440 38048 50456 38112
rect 50520 38048 50536 38112
rect 50600 38048 50608 38112
rect 50288 38047 50608 38048
rect 0 37348 800 37588
rect 4208 37568 4528 37569
rect 4208 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4528 37568
rect 4208 37503 4528 37504
rect 34928 37568 35248 37569
rect 34928 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35248 37568
rect 34928 37503 35248 37504
rect 19568 37024 19888 37025
rect 19568 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19888 37024
rect 19568 36959 19888 36960
rect 50288 37024 50608 37025
rect 50288 36960 50296 37024
rect 50360 36960 50376 37024
rect 50440 36960 50456 37024
rect 50520 36960 50536 37024
rect 50600 36960 50608 37024
rect 50288 36959 50608 36960
rect 59200 36668 60000 36908
rect 4208 36480 4528 36481
rect 4208 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4528 36480
rect 4208 36415 4528 36416
rect 34928 36480 35248 36481
rect 34928 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35248 36480
rect 34928 36415 35248 36416
rect 19568 35936 19888 35937
rect 19568 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19888 35936
rect 19568 35871 19888 35872
rect 50288 35936 50608 35937
rect 50288 35872 50296 35936
rect 50360 35872 50376 35936
rect 50440 35872 50456 35936
rect 50520 35872 50536 35936
rect 50600 35872 50608 35936
rect 50288 35871 50608 35872
rect 4208 35392 4528 35393
rect 4208 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4528 35392
rect 4208 35327 4528 35328
rect 34928 35392 35248 35393
rect 34928 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35248 35392
rect 34928 35327 35248 35328
rect 0 34778 800 34868
rect 19568 34848 19888 34849
rect 19568 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19888 34848
rect 19568 34783 19888 34784
rect 50288 34848 50608 34849
rect 50288 34784 50296 34848
rect 50360 34784 50376 34848
rect 50440 34784 50456 34848
rect 50520 34784 50536 34848
rect 50600 34784 50608 34848
rect 50288 34783 50608 34784
rect 2129 34778 2195 34781
rect 0 34776 2195 34778
rect 0 34720 2134 34776
rect 2190 34720 2195 34776
rect 0 34718 2195 34720
rect 0 34628 800 34718
rect 2129 34715 2195 34718
rect 4208 34304 4528 34305
rect 4208 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4528 34304
rect 4208 34239 4528 34240
rect 34928 34304 35248 34305
rect 34928 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35248 34304
rect 34928 34239 35248 34240
rect 59200 33948 60000 34188
rect 19568 33760 19888 33761
rect 19568 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19888 33760
rect 19568 33695 19888 33696
rect 50288 33760 50608 33761
rect 50288 33696 50296 33760
rect 50360 33696 50376 33760
rect 50440 33696 50456 33760
rect 50520 33696 50536 33760
rect 50600 33696 50608 33760
rect 50288 33695 50608 33696
rect 4208 33216 4528 33217
rect 4208 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4528 33216
rect 4208 33151 4528 33152
rect 34928 33216 35248 33217
rect 34928 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35248 33216
rect 34928 33151 35248 33152
rect 0 32588 800 32828
rect 19568 32672 19888 32673
rect 19568 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19888 32672
rect 19568 32607 19888 32608
rect 50288 32672 50608 32673
rect 50288 32608 50296 32672
rect 50360 32608 50376 32672
rect 50440 32608 50456 32672
rect 50520 32608 50536 32672
rect 50600 32608 50608 32672
rect 50288 32607 50608 32608
rect 4208 32128 4528 32129
rect 4208 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4528 32128
rect 4208 32063 4528 32064
rect 34928 32128 35248 32129
rect 34928 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35248 32128
rect 34928 32063 35248 32064
rect 58157 32058 58223 32061
rect 59200 32058 60000 32148
rect 58157 32056 60000 32058
rect 58157 32000 58162 32056
rect 58218 32000 60000 32056
rect 58157 31998 60000 32000
rect 58157 31995 58223 31998
rect 59200 31908 60000 31998
rect 19568 31584 19888 31585
rect 19568 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19888 31584
rect 19568 31519 19888 31520
rect 50288 31584 50608 31585
rect 50288 31520 50296 31584
rect 50360 31520 50376 31584
rect 50440 31520 50456 31584
rect 50520 31520 50536 31584
rect 50600 31520 50608 31584
rect 50288 31519 50608 31520
rect 4208 31040 4528 31041
rect 4208 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4528 31040
rect 4208 30975 4528 30976
rect 34928 31040 35248 31041
rect 34928 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35248 31040
rect 34928 30975 35248 30976
rect 19568 30496 19888 30497
rect 19568 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19888 30496
rect 19568 30431 19888 30432
rect 50288 30496 50608 30497
rect 50288 30432 50296 30496
rect 50360 30432 50376 30496
rect 50440 30432 50456 30496
rect 50520 30432 50536 30496
rect 50600 30432 50608 30496
rect 50288 30431 50608 30432
rect 0 29868 800 30108
rect 4208 29952 4528 29953
rect 4208 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4528 29952
rect 4208 29887 4528 29888
rect 34928 29952 35248 29953
rect 34928 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35248 29952
rect 34928 29887 35248 29888
rect 19568 29408 19888 29409
rect 19568 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19888 29408
rect 19568 29343 19888 29344
rect 50288 29408 50608 29409
rect 50288 29344 50296 29408
rect 50360 29344 50376 29408
rect 50440 29344 50456 29408
rect 50520 29344 50536 29408
rect 50600 29344 50608 29408
rect 50288 29343 50608 29344
rect 57697 29338 57763 29341
rect 59200 29338 60000 29428
rect 57697 29336 60000 29338
rect 57697 29280 57702 29336
rect 57758 29280 60000 29336
rect 57697 29278 60000 29280
rect 57697 29275 57763 29278
rect 59200 29188 60000 29278
rect 4208 28864 4528 28865
rect 4208 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4528 28864
rect 4208 28799 4528 28800
rect 34928 28864 35248 28865
rect 34928 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35248 28864
rect 34928 28799 35248 28800
rect 19568 28320 19888 28321
rect 19568 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19888 28320
rect 19568 28255 19888 28256
rect 50288 28320 50608 28321
rect 50288 28256 50296 28320
rect 50360 28256 50376 28320
rect 50440 28256 50456 28320
rect 50520 28256 50536 28320
rect 50600 28256 50608 28320
rect 50288 28255 50608 28256
rect 4208 27776 4528 27777
rect 4208 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4528 27776
rect 4208 27711 4528 27712
rect 34928 27776 35248 27777
rect 34928 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35248 27776
rect 34928 27711 35248 27712
rect 0 27148 800 27388
rect 19568 27232 19888 27233
rect 19568 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19888 27232
rect 19568 27167 19888 27168
rect 50288 27232 50608 27233
rect 50288 27168 50296 27232
rect 50360 27168 50376 27232
rect 50440 27168 50456 27232
rect 50520 27168 50536 27232
rect 50600 27168 50608 27232
rect 50288 27167 50608 27168
rect 4208 26688 4528 26689
rect 4208 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4528 26688
rect 4208 26623 4528 26624
rect 34928 26688 35248 26689
rect 34928 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35248 26688
rect 34928 26623 35248 26624
rect 59200 26468 60000 26708
rect 19568 26144 19888 26145
rect 19568 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19888 26144
rect 19568 26079 19888 26080
rect 50288 26144 50608 26145
rect 50288 26080 50296 26144
rect 50360 26080 50376 26144
rect 50440 26080 50456 26144
rect 50520 26080 50536 26144
rect 50600 26080 50608 26144
rect 50288 26079 50608 26080
rect 4208 25600 4528 25601
rect 4208 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4528 25600
rect 4208 25535 4528 25536
rect 34928 25600 35248 25601
rect 34928 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35248 25600
rect 34928 25535 35248 25536
rect 0 25108 800 25348
rect 19568 25056 19888 25057
rect 19568 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19888 25056
rect 19568 24991 19888 24992
rect 50288 25056 50608 25057
rect 50288 24992 50296 25056
rect 50360 24992 50376 25056
rect 50440 24992 50456 25056
rect 50520 24992 50536 25056
rect 50600 24992 50608 25056
rect 50288 24991 50608 24992
rect 58157 24578 58223 24581
rect 59200 24578 60000 24668
rect 58157 24576 60000 24578
rect 58157 24520 58162 24576
rect 58218 24520 60000 24576
rect 58157 24518 60000 24520
rect 58157 24515 58223 24518
rect 4208 24512 4528 24513
rect 4208 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4528 24512
rect 4208 24447 4528 24448
rect 34928 24512 35248 24513
rect 34928 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35248 24512
rect 34928 24447 35248 24448
rect 59200 24428 60000 24518
rect 19568 23968 19888 23969
rect 19568 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19888 23968
rect 19568 23903 19888 23904
rect 50288 23968 50608 23969
rect 50288 23904 50296 23968
rect 50360 23904 50376 23968
rect 50440 23904 50456 23968
rect 50520 23904 50536 23968
rect 50600 23904 50608 23968
rect 50288 23903 50608 23904
rect 4208 23424 4528 23425
rect 4208 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4528 23424
rect 4208 23359 4528 23360
rect 34928 23424 35248 23425
rect 34928 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35248 23424
rect 34928 23359 35248 23360
rect 19568 22880 19888 22881
rect 19568 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19888 22880
rect 19568 22815 19888 22816
rect 50288 22880 50608 22881
rect 50288 22816 50296 22880
rect 50360 22816 50376 22880
rect 50440 22816 50456 22880
rect 50520 22816 50536 22880
rect 50600 22816 50608 22880
rect 50288 22815 50608 22816
rect 0 22388 800 22628
rect 4208 22336 4528 22337
rect 4208 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4528 22336
rect 4208 22271 4528 22272
rect 34928 22336 35248 22337
rect 34928 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35248 22336
rect 34928 22271 35248 22272
rect 19568 21792 19888 21793
rect 19568 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19888 21792
rect 19568 21727 19888 21728
rect 50288 21792 50608 21793
rect 50288 21728 50296 21792
rect 50360 21728 50376 21792
rect 50440 21728 50456 21792
rect 50520 21728 50536 21792
rect 50600 21728 50608 21792
rect 50288 21727 50608 21728
rect 59200 21708 60000 21948
rect 4208 21248 4528 21249
rect 4208 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4528 21248
rect 4208 21183 4528 21184
rect 34928 21248 35248 21249
rect 34928 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35248 21248
rect 34928 21183 35248 21184
rect 19568 20704 19888 20705
rect 19568 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19888 20704
rect 19568 20639 19888 20640
rect 50288 20704 50608 20705
rect 50288 20640 50296 20704
rect 50360 20640 50376 20704
rect 50440 20640 50456 20704
rect 50520 20640 50536 20704
rect 50600 20640 50608 20704
rect 50288 20639 50608 20640
rect 4208 20160 4528 20161
rect 4208 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4528 20160
rect 4208 20095 4528 20096
rect 34928 20160 35248 20161
rect 34928 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35248 20160
rect 34928 20095 35248 20096
rect 0 19668 800 19908
rect 19568 19616 19888 19617
rect 19568 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19888 19616
rect 19568 19551 19888 19552
rect 50288 19616 50608 19617
rect 50288 19552 50296 19616
rect 50360 19552 50376 19616
rect 50440 19552 50456 19616
rect 50520 19552 50536 19616
rect 50600 19552 50608 19616
rect 50288 19551 50608 19552
rect 58157 19138 58223 19141
rect 59200 19138 60000 19228
rect 58157 19136 60000 19138
rect 58157 19080 58162 19136
rect 58218 19080 60000 19136
rect 58157 19078 60000 19080
rect 58157 19075 58223 19078
rect 4208 19072 4528 19073
rect 4208 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4528 19072
rect 4208 19007 4528 19008
rect 34928 19072 35248 19073
rect 34928 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35248 19072
rect 34928 19007 35248 19008
rect 59200 18988 60000 19078
rect 19568 18528 19888 18529
rect 19568 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19888 18528
rect 19568 18463 19888 18464
rect 50288 18528 50608 18529
rect 50288 18464 50296 18528
rect 50360 18464 50376 18528
rect 50440 18464 50456 18528
rect 50520 18464 50536 18528
rect 50600 18464 50608 18528
rect 50288 18463 50608 18464
rect 4208 17984 4528 17985
rect 4208 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4528 17984
rect 4208 17919 4528 17920
rect 34928 17984 35248 17985
rect 34928 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35248 17984
rect 34928 17919 35248 17920
rect 19568 17440 19888 17441
rect 19568 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19888 17440
rect 19568 17375 19888 17376
rect 50288 17440 50608 17441
rect 50288 17376 50296 17440
rect 50360 17376 50376 17440
rect 50440 17376 50456 17440
rect 50520 17376 50536 17440
rect 50600 17376 50608 17440
rect 50288 17375 50608 17376
rect 0 16948 800 17188
rect 4208 16896 4528 16897
rect 4208 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4528 16896
rect 4208 16831 4528 16832
rect 34928 16896 35248 16897
rect 34928 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35248 16896
rect 34928 16831 35248 16832
rect 19568 16352 19888 16353
rect 19568 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19888 16352
rect 19568 16287 19888 16288
rect 50288 16352 50608 16353
rect 50288 16288 50296 16352
rect 50360 16288 50376 16352
rect 50440 16288 50456 16352
rect 50520 16288 50536 16352
rect 50600 16288 50608 16352
rect 50288 16287 50608 16288
rect 59200 16268 60000 16508
rect 4208 15808 4528 15809
rect 4208 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4528 15808
rect 4208 15743 4528 15744
rect 34928 15808 35248 15809
rect 34928 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35248 15808
rect 34928 15743 35248 15744
rect 19568 15264 19888 15265
rect 19568 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19888 15264
rect 19568 15199 19888 15200
rect 50288 15264 50608 15265
rect 50288 15200 50296 15264
rect 50360 15200 50376 15264
rect 50440 15200 50456 15264
rect 50520 15200 50536 15264
rect 50600 15200 50608 15264
rect 50288 15199 50608 15200
rect 0 14908 800 15148
rect 4208 14720 4528 14721
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 4208 14655 4528 14656
rect 34928 14720 35248 14721
rect 34928 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35248 14720
rect 34928 14655 35248 14656
rect 59200 14228 60000 14468
rect 19568 14176 19888 14177
rect 19568 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19888 14176
rect 19568 14111 19888 14112
rect 50288 14176 50608 14177
rect 50288 14112 50296 14176
rect 50360 14112 50376 14176
rect 50440 14112 50456 14176
rect 50520 14112 50536 14176
rect 50600 14112 50608 14176
rect 50288 14111 50608 14112
rect 4208 13632 4528 13633
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 13567 4528 13568
rect 34928 13632 35248 13633
rect 34928 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35248 13632
rect 34928 13567 35248 13568
rect 19568 13088 19888 13089
rect 19568 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19888 13088
rect 19568 13023 19888 13024
rect 50288 13088 50608 13089
rect 50288 13024 50296 13088
rect 50360 13024 50376 13088
rect 50440 13024 50456 13088
rect 50520 13024 50536 13088
rect 50600 13024 50608 13088
rect 50288 13023 50608 13024
rect 4208 12544 4528 12545
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 12479 4528 12480
rect 34928 12544 35248 12545
rect 34928 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35248 12544
rect 34928 12479 35248 12480
rect 0 12188 800 12428
rect 19568 12000 19888 12001
rect 19568 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19888 12000
rect 19568 11935 19888 11936
rect 50288 12000 50608 12001
rect 50288 11936 50296 12000
rect 50360 11936 50376 12000
rect 50440 11936 50456 12000
rect 50520 11936 50536 12000
rect 50600 11936 50608 12000
rect 50288 11935 50608 11936
rect 58157 11658 58223 11661
rect 59200 11658 60000 11748
rect 58157 11656 60000 11658
rect 58157 11600 58162 11656
rect 58218 11600 60000 11656
rect 58157 11598 60000 11600
rect 58157 11595 58223 11598
rect 59200 11508 60000 11598
rect 4208 11456 4528 11457
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 11391 4528 11392
rect 34928 11456 35248 11457
rect 34928 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35248 11456
rect 34928 11391 35248 11392
rect 19568 10912 19888 10913
rect 19568 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19888 10912
rect 19568 10847 19888 10848
rect 50288 10912 50608 10913
rect 50288 10848 50296 10912
rect 50360 10848 50376 10912
rect 50440 10848 50456 10912
rect 50520 10848 50536 10912
rect 50600 10848 50608 10912
rect 50288 10847 50608 10848
rect 4208 10368 4528 10369
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 10303 4528 10304
rect 34928 10368 35248 10369
rect 34928 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35248 10368
rect 34928 10303 35248 10304
rect 19568 9824 19888 9825
rect 19568 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19888 9824
rect 19568 9759 19888 9760
rect 50288 9824 50608 9825
rect 50288 9760 50296 9824
rect 50360 9760 50376 9824
rect 50440 9760 50456 9824
rect 50520 9760 50536 9824
rect 50600 9760 50608 9824
rect 50288 9759 50608 9760
rect 0 9618 800 9708
rect 2773 9618 2839 9621
rect 0 9616 2839 9618
rect 0 9560 2778 9616
rect 2834 9560 2839 9616
rect 0 9558 2839 9560
rect 0 9468 800 9558
rect 2773 9555 2839 9558
rect 4208 9280 4528 9281
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 9215 4528 9216
rect 34928 9280 35248 9281
rect 34928 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35248 9280
rect 34928 9215 35248 9216
rect 58157 8938 58223 8941
rect 59200 8938 60000 9028
rect 58157 8936 60000 8938
rect 58157 8880 58162 8936
rect 58218 8880 60000 8936
rect 58157 8878 60000 8880
rect 58157 8875 58223 8878
rect 59200 8788 60000 8878
rect 19568 8736 19888 8737
rect 19568 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19888 8736
rect 19568 8671 19888 8672
rect 50288 8736 50608 8737
rect 50288 8672 50296 8736
rect 50360 8672 50376 8736
rect 50440 8672 50456 8736
rect 50520 8672 50536 8736
rect 50600 8672 50608 8736
rect 50288 8671 50608 8672
rect 4208 8192 4528 8193
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 8127 4528 8128
rect 34928 8192 35248 8193
rect 34928 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35248 8192
rect 34928 8127 35248 8128
rect 0 7428 800 7668
rect 19568 7648 19888 7649
rect 19568 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19888 7648
rect 19568 7583 19888 7584
rect 50288 7648 50608 7649
rect 50288 7584 50296 7648
rect 50360 7584 50376 7648
rect 50440 7584 50456 7648
rect 50520 7584 50536 7648
rect 50600 7584 50608 7648
rect 50288 7583 50608 7584
rect 4208 7104 4528 7105
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 7039 4528 7040
rect 34928 7104 35248 7105
rect 34928 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35248 7104
rect 34928 7039 35248 7040
rect 59200 6748 60000 6988
rect 19568 6560 19888 6561
rect 19568 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19888 6560
rect 19568 6495 19888 6496
rect 50288 6560 50608 6561
rect 50288 6496 50296 6560
rect 50360 6496 50376 6560
rect 50440 6496 50456 6560
rect 50520 6496 50536 6560
rect 50600 6496 50608 6560
rect 50288 6495 50608 6496
rect 4208 6016 4528 6017
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 5951 4528 5952
rect 34928 6016 35248 6017
rect 34928 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35248 6016
rect 34928 5951 35248 5952
rect 19568 5472 19888 5473
rect 19568 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19888 5472
rect 19568 5407 19888 5408
rect 50288 5472 50608 5473
rect 50288 5408 50296 5472
rect 50360 5408 50376 5472
rect 50440 5408 50456 5472
rect 50520 5408 50536 5472
rect 50600 5408 50608 5472
rect 50288 5407 50608 5408
rect 0 4858 800 4948
rect 4208 4928 4528 4929
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 4863 4528 4864
rect 34928 4928 35248 4929
rect 34928 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35248 4928
rect 34928 4863 35248 4864
rect 2773 4858 2839 4861
rect 0 4856 2839 4858
rect 0 4800 2778 4856
rect 2834 4800 2839 4856
rect 0 4798 2839 4800
rect 0 4708 800 4798
rect 2773 4795 2839 4798
rect 19568 4384 19888 4385
rect 19568 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19888 4384
rect 19568 4319 19888 4320
rect 50288 4384 50608 4385
rect 50288 4320 50296 4384
rect 50360 4320 50376 4384
rect 50440 4320 50456 4384
rect 50520 4320 50536 4384
rect 50600 4320 50608 4384
rect 50288 4319 50608 4320
rect 59200 4028 60000 4268
rect 4208 3840 4528 3841
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 3775 4528 3776
rect 34928 3840 35248 3841
rect 34928 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35248 3840
rect 34928 3775 35248 3776
rect 19568 3296 19888 3297
rect 19568 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19888 3296
rect 19568 3231 19888 3232
rect 50288 3296 50608 3297
rect 50288 3232 50296 3296
rect 50360 3232 50376 3296
rect 50440 3232 50456 3296
rect 50520 3232 50536 3296
rect 50600 3232 50608 3296
rect 50288 3231 50608 3232
rect 4208 2752 4528 2753
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2687 4528 2688
rect 34928 2752 35248 2753
rect 34928 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35248 2752
rect 34928 2687 35248 2688
rect 0 1988 800 2228
rect 19568 2208 19888 2209
rect 19568 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19888 2208
rect 19568 2143 19888 2144
rect 50288 2208 50608 2209
rect 50288 2144 50296 2208
rect 50360 2144 50376 2208
rect 50440 2144 50456 2208
rect 50520 2144 50536 2208
rect 50600 2144 50608 2208
rect 50288 2143 50608 2144
rect 57881 1458 57947 1461
rect 59200 1458 60000 1548
rect 57881 1456 60000 1458
rect 57881 1400 57886 1456
rect 57942 1400 60000 1456
rect 57881 1398 60000 1400
rect 57881 1395 57947 1398
rect 59200 1308 60000 1398
<< via3 >>
rect 19576 57692 19640 57696
rect 19576 57636 19580 57692
rect 19580 57636 19636 57692
rect 19636 57636 19640 57692
rect 19576 57632 19640 57636
rect 19656 57692 19720 57696
rect 19656 57636 19660 57692
rect 19660 57636 19716 57692
rect 19716 57636 19720 57692
rect 19656 57632 19720 57636
rect 19736 57692 19800 57696
rect 19736 57636 19740 57692
rect 19740 57636 19796 57692
rect 19796 57636 19800 57692
rect 19736 57632 19800 57636
rect 19816 57692 19880 57696
rect 19816 57636 19820 57692
rect 19820 57636 19876 57692
rect 19876 57636 19880 57692
rect 19816 57632 19880 57636
rect 50296 57692 50360 57696
rect 50296 57636 50300 57692
rect 50300 57636 50356 57692
rect 50356 57636 50360 57692
rect 50296 57632 50360 57636
rect 50376 57692 50440 57696
rect 50376 57636 50380 57692
rect 50380 57636 50436 57692
rect 50436 57636 50440 57692
rect 50376 57632 50440 57636
rect 50456 57692 50520 57696
rect 50456 57636 50460 57692
rect 50460 57636 50516 57692
rect 50516 57636 50520 57692
rect 50456 57632 50520 57636
rect 50536 57692 50600 57696
rect 50536 57636 50540 57692
rect 50540 57636 50596 57692
rect 50596 57636 50600 57692
rect 50536 57632 50600 57636
rect 4216 57148 4280 57152
rect 4216 57092 4220 57148
rect 4220 57092 4276 57148
rect 4276 57092 4280 57148
rect 4216 57088 4280 57092
rect 4296 57148 4360 57152
rect 4296 57092 4300 57148
rect 4300 57092 4356 57148
rect 4356 57092 4360 57148
rect 4296 57088 4360 57092
rect 4376 57148 4440 57152
rect 4376 57092 4380 57148
rect 4380 57092 4436 57148
rect 4436 57092 4440 57148
rect 4376 57088 4440 57092
rect 4456 57148 4520 57152
rect 4456 57092 4460 57148
rect 4460 57092 4516 57148
rect 4516 57092 4520 57148
rect 4456 57088 4520 57092
rect 34936 57148 35000 57152
rect 34936 57092 34940 57148
rect 34940 57092 34996 57148
rect 34996 57092 35000 57148
rect 34936 57088 35000 57092
rect 35016 57148 35080 57152
rect 35016 57092 35020 57148
rect 35020 57092 35076 57148
rect 35076 57092 35080 57148
rect 35016 57088 35080 57092
rect 35096 57148 35160 57152
rect 35096 57092 35100 57148
rect 35100 57092 35156 57148
rect 35156 57092 35160 57148
rect 35096 57088 35160 57092
rect 35176 57148 35240 57152
rect 35176 57092 35180 57148
rect 35180 57092 35236 57148
rect 35236 57092 35240 57148
rect 35176 57088 35240 57092
rect 19576 56604 19640 56608
rect 19576 56548 19580 56604
rect 19580 56548 19636 56604
rect 19636 56548 19640 56604
rect 19576 56544 19640 56548
rect 19656 56604 19720 56608
rect 19656 56548 19660 56604
rect 19660 56548 19716 56604
rect 19716 56548 19720 56604
rect 19656 56544 19720 56548
rect 19736 56604 19800 56608
rect 19736 56548 19740 56604
rect 19740 56548 19796 56604
rect 19796 56548 19800 56604
rect 19736 56544 19800 56548
rect 19816 56604 19880 56608
rect 19816 56548 19820 56604
rect 19820 56548 19876 56604
rect 19876 56548 19880 56604
rect 19816 56544 19880 56548
rect 50296 56604 50360 56608
rect 50296 56548 50300 56604
rect 50300 56548 50356 56604
rect 50356 56548 50360 56604
rect 50296 56544 50360 56548
rect 50376 56604 50440 56608
rect 50376 56548 50380 56604
rect 50380 56548 50436 56604
rect 50436 56548 50440 56604
rect 50376 56544 50440 56548
rect 50456 56604 50520 56608
rect 50456 56548 50460 56604
rect 50460 56548 50516 56604
rect 50516 56548 50520 56604
rect 50456 56544 50520 56548
rect 50536 56604 50600 56608
rect 50536 56548 50540 56604
rect 50540 56548 50596 56604
rect 50596 56548 50600 56604
rect 50536 56544 50600 56548
rect 4216 56060 4280 56064
rect 4216 56004 4220 56060
rect 4220 56004 4276 56060
rect 4276 56004 4280 56060
rect 4216 56000 4280 56004
rect 4296 56060 4360 56064
rect 4296 56004 4300 56060
rect 4300 56004 4356 56060
rect 4356 56004 4360 56060
rect 4296 56000 4360 56004
rect 4376 56060 4440 56064
rect 4376 56004 4380 56060
rect 4380 56004 4436 56060
rect 4436 56004 4440 56060
rect 4376 56000 4440 56004
rect 4456 56060 4520 56064
rect 4456 56004 4460 56060
rect 4460 56004 4516 56060
rect 4516 56004 4520 56060
rect 4456 56000 4520 56004
rect 34936 56060 35000 56064
rect 34936 56004 34940 56060
rect 34940 56004 34996 56060
rect 34996 56004 35000 56060
rect 34936 56000 35000 56004
rect 35016 56060 35080 56064
rect 35016 56004 35020 56060
rect 35020 56004 35076 56060
rect 35076 56004 35080 56060
rect 35016 56000 35080 56004
rect 35096 56060 35160 56064
rect 35096 56004 35100 56060
rect 35100 56004 35156 56060
rect 35156 56004 35160 56060
rect 35096 56000 35160 56004
rect 35176 56060 35240 56064
rect 35176 56004 35180 56060
rect 35180 56004 35236 56060
rect 35236 56004 35240 56060
rect 35176 56000 35240 56004
rect 19576 55516 19640 55520
rect 19576 55460 19580 55516
rect 19580 55460 19636 55516
rect 19636 55460 19640 55516
rect 19576 55456 19640 55460
rect 19656 55516 19720 55520
rect 19656 55460 19660 55516
rect 19660 55460 19716 55516
rect 19716 55460 19720 55516
rect 19656 55456 19720 55460
rect 19736 55516 19800 55520
rect 19736 55460 19740 55516
rect 19740 55460 19796 55516
rect 19796 55460 19800 55516
rect 19736 55456 19800 55460
rect 19816 55516 19880 55520
rect 19816 55460 19820 55516
rect 19820 55460 19876 55516
rect 19876 55460 19880 55516
rect 19816 55456 19880 55460
rect 50296 55516 50360 55520
rect 50296 55460 50300 55516
rect 50300 55460 50356 55516
rect 50356 55460 50360 55516
rect 50296 55456 50360 55460
rect 50376 55516 50440 55520
rect 50376 55460 50380 55516
rect 50380 55460 50436 55516
rect 50436 55460 50440 55516
rect 50376 55456 50440 55460
rect 50456 55516 50520 55520
rect 50456 55460 50460 55516
rect 50460 55460 50516 55516
rect 50516 55460 50520 55516
rect 50456 55456 50520 55460
rect 50536 55516 50600 55520
rect 50536 55460 50540 55516
rect 50540 55460 50596 55516
rect 50596 55460 50600 55516
rect 50536 55456 50600 55460
rect 4216 54972 4280 54976
rect 4216 54916 4220 54972
rect 4220 54916 4276 54972
rect 4276 54916 4280 54972
rect 4216 54912 4280 54916
rect 4296 54972 4360 54976
rect 4296 54916 4300 54972
rect 4300 54916 4356 54972
rect 4356 54916 4360 54972
rect 4296 54912 4360 54916
rect 4376 54972 4440 54976
rect 4376 54916 4380 54972
rect 4380 54916 4436 54972
rect 4436 54916 4440 54972
rect 4376 54912 4440 54916
rect 4456 54972 4520 54976
rect 4456 54916 4460 54972
rect 4460 54916 4516 54972
rect 4516 54916 4520 54972
rect 4456 54912 4520 54916
rect 34936 54972 35000 54976
rect 34936 54916 34940 54972
rect 34940 54916 34996 54972
rect 34996 54916 35000 54972
rect 34936 54912 35000 54916
rect 35016 54972 35080 54976
rect 35016 54916 35020 54972
rect 35020 54916 35076 54972
rect 35076 54916 35080 54972
rect 35016 54912 35080 54916
rect 35096 54972 35160 54976
rect 35096 54916 35100 54972
rect 35100 54916 35156 54972
rect 35156 54916 35160 54972
rect 35096 54912 35160 54916
rect 35176 54972 35240 54976
rect 35176 54916 35180 54972
rect 35180 54916 35236 54972
rect 35236 54916 35240 54972
rect 35176 54912 35240 54916
rect 19576 54428 19640 54432
rect 19576 54372 19580 54428
rect 19580 54372 19636 54428
rect 19636 54372 19640 54428
rect 19576 54368 19640 54372
rect 19656 54428 19720 54432
rect 19656 54372 19660 54428
rect 19660 54372 19716 54428
rect 19716 54372 19720 54428
rect 19656 54368 19720 54372
rect 19736 54428 19800 54432
rect 19736 54372 19740 54428
rect 19740 54372 19796 54428
rect 19796 54372 19800 54428
rect 19736 54368 19800 54372
rect 19816 54428 19880 54432
rect 19816 54372 19820 54428
rect 19820 54372 19876 54428
rect 19876 54372 19880 54428
rect 19816 54368 19880 54372
rect 50296 54428 50360 54432
rect 50296 54372 50300 54428
rect 50300 54372 50356 54428
rect 50356 54372 50360 54428
rect 50296 54368 50360 54372
rect 50376 54428 50440 54432
rect 50376 54372 50380 54428
rect 50380 54372 50436 54428
rect 50436 54372 50440 54428
rect 50376 54368 50440 54372
rect 50456 54428 50520 54432
rect 50456 54372 50460 54428
rect 50460 54372 50516 54428
rect 50516 54372 50520 54428
rect 50456 54368 50520 54372
rect 50536 54428 50600 54432
rect 50536 54372 50540 54428
rect 50540 54372 50596 54428
rect 50596 54372 50600 54428
rect 50536 54368 50600 54372
rect 4216 53884 4280 53888
rect 4216 53828 4220 53884
rect 4220 53828 4276 53884
rect 4276 53828 4280 53884
rect 4216 53824 4280 53828
rect 4296 53884 4360 53888
rect 4296 53828 4300 53884
rect 4300 53828 4356 53884
rect 4356 53828 4360 53884
rect 4296 53824 4360 53828
rect 4376 53884 4440 53888
rect 4376 53828 4380 53884
rect 4380 53828 4436 53884
rect 4436 53828 4440 53884
rect 4376 53824 4440 53828
rect 4456 53884 4520 53888
rect 4456 53828 4460 53884
rect 4460 53828 4516 53884
rect 4516 53828 4520 53884
rect 4456 53824 4520 53828
rect 34936 53884 35000 53888
rect 34936 53828 34940 53884
rect 34940 53828 34996 53884
rect 34996 53828 35000 53884
rect 34936 53824 35000 53828
rect 35016 53884 35080 53888
rect 35016 53828 35020 53884
rect 35020 53828 35076 53884
rect 35076 53828 35080 53884
rect 35016 53824 35080 53828
rect 35096 53884 35160 53888
rect 35096 53828 35100 53884
rect 35100 53828 35156 53884
rect 35156 53828 35160 53884
rect 35096 53824 35160 53828
rect 35176 53884 35240 53888
rect 35176 53828 35180 53884
rect 35180 53828 35236 53884
rect 35236 53828 35240 53884
rect 35176 53824 35240 53828
rect 19576 53340 19640 53344
rect 19576 53284 19580 53340
rect 19580 53284 19636 53340
rect 19636 53284 19640 53340
rect 19576 53280 19640 53284
rect 19656 53340 19720 53344
rect 19656 53284 19660 53340
rect 19660 53284 19716 53340
rect 19716 53284 19720 53340
rect 19656 53280 19720 53284
rect 19736 53340 19800 53344
rect 19736 53284 19740 53340
rect 19740 53284 19796 53340
rect 19796 53284 19800 53340
rect 19736 53280 19800 53284
rect 19816 53340 19880 53344
rect 19816 53284 19820 53340
rect 19820 53284 19876 53340
rect 19876 53284 19880 53340
rect 19816 53280 19880 53284
rect 50296 53340 50360 53344
rect 50296 53284 50300 53340
rect 50300 53284 50356 53340
rect 50356 53284 50360 53340
rect 50296 53280 50360 53284
rect 50376 53340 50440 53344
rect 50376 53284 50380 53340
rect 50380 53284 50436 53340
rect 50436 53284 50440 53340
rect 50376 53280 50440 53284
rect 50456 53340 50520 53344
rect 50456 53284 50460 53340
rect 50460 53284 50516 53340
rect 50516 53284 50520 53340
rect 50456 53280 50520 53284
rect 50536 53340 50600 53344
rect 50536 53284 50540 53340
rect 50540 53284 50596 53340
rect 50596 53284 50600 53340
rect 50536 53280 50600 53284
rect 4216 52796 4280 52800
rect 4216 52740 4220 52796
rect 4220 52740 4276 52796
rect 4276 52740 4280 52796
rect 4216 52736 4280 52740
rect 4296 52796 4360 52800
rect 4296 52740 4300 52796
rect 4300 52740 4356 52796
rect 4356 52740 4360 52796
rect 4296 52736 4360 52740
rect 4376 52796 4440 52800
rect 4376 52740 4380 52796
rect 4380 52740 4436 52796
rect 4436 52740 4440 52796
rect 4376 52736 4440 52740
rect 4456 52796 4520 52800
rect 4456 52740 4460 52796
rect 4460 52740 4516 52796
rect 4516 52740 4520 52796
rect 4456 52736 4520 52740
rect 34936 52796 35000 52800
rect 34936 52740 34940 52796
rect 34940 52740 34996 52796
rect 34996 52740 35000 52796
rect 34936 52736 35000 52740
rect 35016 52796 35080 52800
rect 35016 52740 35020 52796
rect 35020 52740 35076 52796
rect 35076 52740 35080 52796
rect 35016 52736 35080 52740
rect 35096 52796 35160 52800
rect 35096 52740 35100 52796
rect 35100 52740 35156 52796
rect 35156 52740 35160 52796
rect 35096 52736 35160 52740
rect 35176 52796 35240 52800
rect 35176 52740 35180 52796
rect 35180 52740 35236 52796
rect 35236 52740 35240 52796
rect 35176 52736 35240 52740
rect 19576 52252 19640 52256
rect 19576 52196 19580 52252
rect 19580 52196 19636 52252
rect 19636 52196 19640 52252
rect 19576 52192 19640 52196
rect 19656 52252 19720 52256
rect 19656 52196 19660 52252
rect 19660 52196 19716 52252
rect 19716 52196 19720 52252
rect 19656 52192 19720 52196
rect 19736 52252 19800 52256
rect 19736 52196 19740 52252
rect 19740 52196 19796 52252
rect 19796 52196 19800 52252
rect 19736 52192 19800 52196
rect 19816 52252 19880 52256
rect 19816 52196 19820 52252
rect 19820 52196 19876 52252
rect 19876 52196 19880 52252
rect 19816 52192 19880 52196
rect 50296 52252 50360 52256
rect 50296 52196 50300 52252
rect 50300 52196 50356 52252
rect 50356 52196 50360 52252
rect 50296 52192 50360 52196
rect 50376 52252 50440 52256
rect 50376 52196 50380 52252
rect 50380 52196 50436 52252
rect 50436 52196 50440 52252
rect 50376 52192 50440 52196
rect 50456 52252 50520 52256
rect 50456 52196 50460 52252
rect 50460 52196 50516 52252
rect 50516 52196 50520 52252
rect 50456 52192 50520 52196
rect 50536 52252 50600 52256
rect 50536 52196 50540 52252
rect 50540 52196 50596 52252
rect 50596 52196 50600 52252
rect 50536 52192 50600 52196
rect 4216 51708 4280 51712
rect 4216 51652 4220 51708
rect 4220 51652 4276 51708
rect 4276 51652 4280 51708
rect 4216 51648 4280 51652
rect 4296 51708 4360 51712
rect 4296 51652 4300 51708
rect 4300 51652 4356 51708
rect 4356 51652 4360 51708
rect 4296 51648 4360 51652
rect 4376 51708 4440 51712
rect 4376 51652 4380 51708
rect 4380 51652 4436 51708
rect 4436 51652 4440 51708
rect 4376 51648 4440 51652
rect 4456 51708 4520 51712
rect 4456 51652 4460 51708
rect 4460 51652 4516 51708
rect 4516 51652 4520 51708
rect 4456 51648 4520 51652
rect 34936 51708 35000 51712
rect 34936 51652 34940 51708
rect 34940 51652 34996 51708
rect 34996 51652 35000 51708
rect 34936 51648 35000 51652
rect 35016 51708 35080 51712
rect 35016 51652 35020 51708
rect 35020 51652 35076 51708
rect 35076 51652 35080 51708
rect 35016 51648 35080 51652
rect 35096 51708 35160 51712
rect 35096 51652 35100 51708
rect 35100 51652 35156 51708
rect 35156 51652 35160 51708
rect 35096 51648 35160 51652
rect 35176 51708 35240 51712
rect 35176 51652 35180 51708
rect 35180 51652 35236 51708
rect 35236 51652 35240 51708
rect 35176 51648 35240 51652
rect 19576 51164 19640 51168
rect 19576 51108 19580 51164
rect 19580 51108 19636 51164
rect 19636 51108 19640 51164
rect 19576 51104 19640 51108
rect 19656 51164 19720 51168
rect 19656 51108 19660 51164
rect 19660 51108 19716 51164
rect 19716 51108 19720 51164
rect 19656 51104 19720 51108
rect 19736 51164 19800 51168
rect 19736 51108 19740 51164
rect 19740 51108 19796 51164
rect 19796 51108 19800 51164
rect 19736 51104 19800 51108
rect 19816 51164 19880 51168
rect 19816 51108 19820 51164
rect 19820 51108 19876 51164
rect 19876 51108 19880 51164
rect 19816 51104 19880 51108
rect 50296 51164 50360 51168
rect 50296 51108 50300 51164
rect 50300 51108 50356 51164
rect 50356 51108 50360 51164
rect 50296 51104 50360 51108
rect 50376 51164 50440 51168
rect 50376 51108 50380 51164
rect 50380 51108 50436 51164
rect 50436 51108 50440 51164
rect 50376 51104 50440 51108
rect 50456 51164 50520 51168
rect 50456 51108 50460 51164
rect 50460 51108 50516 51164
rect 50516 51108 50520 51164
rect 50456 51104 50520 51108
rect 50536 51164 50600 51168
rect 50536 51108 50540 51164
rect 50540 51108 50596 51164
rect 50596 51108 50600 51164
rect 50536 51104 50600 51108
rect 4216 50620 4280 50624
rect 4216 50564 4220 50620
rect 4220 50564 4276 50620
rect 4276 50564 4280 50620
rect 4216 50560 4280 50564
rect 4296 50620 4360 50624
rect 4296 50564 4300 50620
rect 4300 50564 4356 50620
rect 4356 50564 4360 50620
rect 4296 50560 4360 50564
rect 4376 50620 4440 50624
rect 4376 50564 4380 50620
rect 4380 50564 4436 50620
rect 4436 50564 4440 50620
rect 4376 50560 4440 50564
rect 4456 50620 4520 50624
rect 4456 50564 4460 50620
rect 4460 50564 4516 50620
rect 4516 50564 4520 50620
rect 4456 50560 4520 50564
rect 34936 50620 35000 50624
rect 34936 50564 34940 50620
rect 34940 50564 34996 50620
rect 34996 50564 35000 50620
rect 34936 50560 35000 50564
rect 35016 50620 35080 50624
rect 35016 50564 35020 50620
rect 35020 50564 35076 50620
rect 35076 50564 35080 50620
rect 35016 50560 35080 50564
rect 35096 50620 35160 50624
rect 35096 50564 35100 50620
rect 35100 50564 35156 50620
rect 35156 50564 35160 50620
rect 35096 50560 35160 50564
rect 35176 50620 35240 50624
rect 35176 50564 35180 50620
rect 35180 50564 35236 50620
rect 35236 50564 35240 50620
rect 35176 50560 35240 50564
rect 19576 50076 19640 50080
rect 19576 50020 19580 50076
rect 19580 50020 19636 50076
rect 19636 50020 19640 50076
rect 19576 50016 19640 50020
rect 19656 50076 19720 50080
rect 19656 50020 19660 50076
rect 19660 50020 19716 50076
rect 19716 50020 19720 50076
rect 19656 50016 19720 50020
rect 19736 50076 19800 50080
rect 19736 50020 19740 50076
rect 19740 50020 19796 50076
rect 19796 50020 19800 50076
rect 19736 50016 19800 50020
rect 19816 50076 19880 50080
rect 19816 50020 19820 50076
rect 19820 50020 19876 50076
rect 19876 50020 19880 50076
rect 19816 50016 19880 50020
rect 50296 50076 50360 50080
rect 50296 50020 50300 50076
rect 50300 50020 50356 50076
rect 50356 50020 50360 50076
rect 50296 50016 50360 50020
rect 50376 50076 50440 50080
rect 50376 50020 50380 50076
rect 50380 50020 50436 50076
rect 50436 50020 50440 50076
rect 50376 50016 50440 50020
rect 50456 50076 50520 50080
rect 50456 50020 50460 50076
rect 50460 50020 50516 50076
rect 50516 50020 50520 50076
rect 50456 50016 50520 50020
rect 50536 50076 50600 50080
rect 50536 50020 50540 50076
rect 50540 50020 50596 50076
rect 50596 50020 50600 50076
rect 50536 50016 50600 50020
rect 4216 49532 4280 49536
rect 4216 49476 4220 49532
rect 4220 49476 4276 49532
rect 4276 49476 4280 49532
rect 4216 49472 4280 49476
rect 4296 49532 4360 49536
rect 4296 49476 4300 49532
rect 4300 49476 4356 49532
rect 4356 49476 4360 49532
rect 4296 49472 4360 49476
rect 4376 49532 4440 49536
rect 4376 49476 4380 49532
rect 4380 49476 4436 49532
rect 4436 49476 4440 49532
rect 4376 49472 4440 49476
rect 4456 49532 4520 49536
rect 4456 49476 4460 49532
rect 4460 49476 4516 49532
rect 4516 49476 4520 49532
rect 4456 49472 4520 49476
rect 34936 49532 35000 49536
rect 34936 49476 34940 49532
rect 34940 49476 34996 49532
rect 34996 49476 35000 49532
rect 34936 49472 35000 49476
rect 35016 49532 35080 49536
rect 35016 49476 35020 49532
rect 35020 49476 35076 49532
rect 35076 49476 35080 49532
rect 35016 49472 35080 49476
rect 35096 49532 35160 49536
rect 35096 49476 35100 49532
rect 35100 49476 35156 49532
rect 35156 49476 35160 49532
rect 35096 49472 35160 49476
rect 35176 49532 35240 49536
rect 35176 49476 35180 49532
rect 35180 49476 35236 49532
rect 35236 49476 35240 49532
rect 35176 49472 35240 49476
rect 19576 48988 19640 48992
rect 19576 48932 19580 48988
rect 19580 48932 19636 48988
rect 19636 48932 19640 48988
rect 19576 48928 19640 48932
rect 19656 48988 19720 48992
rect 19656 48932 19660 48988
rect 19660 48932 19716 48988
rect 19716 48932 19720 48988
rect 19656 48928 19720 48932
rect 19736 48988 19800 48992
rect 19736 48932 19740 48988
rect 19740 48932 19796 48988
rect 19796 48932 19800 48988
rect 19736 48928 19800 48932
rect 19816 48988 19880 48992
rect 19816 48932 19820 48988
rect 19820 48932 19876 48988
rect 19876 48932 19880 48988
rect 19816 48928 19880 48932
rect 50296 48988 50360 48992
rect 50296 48932 50300 48988
rect 50300 48932 50356 48988
rect 50356 48932 50360 48988
rect 50296 48928 50360 48932
rect 50376 48988 50440 48992
rect 50376 48932 50380 48988
rect 50380 48932 50436 48988
rect 50436 48932 50440 48988
rect 50376 48928 50440 48932
rect 50456 48988 50520 48992
rect 50456 48932 50460 48988
rect 50460 48932 50516 48988
rect 50516 48932 50520 48988
rect 50456 48928 50520 48932
rect 50536 48988 50600 48992
rect 50536 48932 50540 48988
rect 50540 48932 50596 48988
rect 50596 48932 50600 48988
rect 50536 48928 50600 48932
rect 4216 48444 4280 48448
rect 4216 48388 4220 48444
rect 4220 48388 4276 48444
rect 4276 48388 4280 48444
rect 4216 48384 4280 48388
rect 4296 48444 4360 48448
rect 4296 48388 4300 48444
rect 4300 48388 4356 48444
rect 4356 48388 4360 48444
rect 4296 48384 4360 48388
rect 4376 48444 4440 48448
rect 4376 48388 4380 48444
rect 4380 48388 4436 48444
rect 4436 48388 4440 48444
rect 4376 48384 4440 48388
rect 4456 48444 4520 48448
rect 4456 48388 4460 48444
rect 4460 48388 4516 48444
rect 4516 48388 4520 48444
rect 4456 48384 4520 48388
rect 34936 48444 35000 48448
rect 34936 48388 34940 48444
rect 34940 48388 34996 48444
rect 34996 48388 35000 48444
rect 34936 48384 35000 48388
rect 35016 48444 35080 48448
rect 35016 48388 35020 48444
rect 35020 48388 35076 48444
rect 35076 48388 35080 48444
rect 35016 48384 35080 48388
rect 35096 48444 35160 48448
rect 35096 48388 35100 48444
rect 35100 48388 35156 48444
rect 35156 48388 35160 48444
rect 35096 48384 35160 48388
rect 35176 48444 35240 48448
rect 35176 48388 35180 48444
rect 35180 48388 35236 48444
rect 35236 48388 35240 48444
rect 35176 48384 35240 48388
rect 19576 47900 19640 47904
rect 19576 47844 19580 47900
rect 19580 47844 19636 47900
rect 19636 47844 19640 47900
rect 19576 47840 19640 47844
rect 19656 47900 19720 47904
rect 19656 47844 19660 47900
rect 19660 47844 19716 47900
rect 19716 47844 19720 47900
rect 19656 47840 19720 47844
rect 19736 47900 19800 47904
rect 19736 47844 19740 47900
rect 19740 47844 19796 47900
rect 19796 47844 19800 47900
rect 19736 47840 19800 47844
rect 19816 47900 19880 47904
rect 19816 47844 19820 47900
rect 19820 47844 19876 47900
rect 19876 47844 19880 47900
rect 19816 47840 19880 47844
rect 50296 47900 50360 47904
rect 50296 47844 50300 47900
rect 50300 47844 50356 47900
rect 50356 47844 50360 47900
rect 50296 47840 50360 47844
rect 50376 47900 50440 47904
rect 50376 47844 50380 47900
rect 50380 47844 50436 47900
rect 50436 47844 50440 47900
rect 50376 47840 50440 47844
rect 50456 47900 50520 47904
rect 50456 47844 50460 47900
rect 50460 47844 50516 47900
rect 50516 47844 50520 47900
rect 50456 47840 50520 47844
rect 50536 47900 50600 47904
rect 50536 47844 50540 47900
rect 50540 47844 50596 47900
rect 50596 47844 50600 47900
rect 50536 47840 50600 47844
rect 4216 47356 4280 47360
rect 4216 47300 4220 47356
rect 4220 47300 4276 47356
rect 4276 47300 4280 47356
rect 4216 47296 4280 47300
rect 4296 47356 4360 47360
rect 4296 47300 4300 47356
rect 4300 47300 4356 47356
rect 4356 47300 4360 47356
rect 4296 47296 4360 47300
rect 4376 47356 4440 47360
rect 4376 47300 4380 47356
rect 4380 47300 4436 47356
rect 4436 47300 4440 47356
rect 4376 47296 4440 47300
rect 4456 47356 4520 47360
rect 4456 47300 4460 47356
rect 4460 47300 4516 47356
rect 4516 47300 4520 47356
rect 4456 47296 4520 47300
rect 34936 47356 35000 47360
rect 34936 47300 34940 47356
rect 34940 47300 34996 47356
rect 34996 47300 35000 47356
rect 34936 47296 35000 47300
rect 35016 47356 35080 47360
rect 35016 47300 35020 47356
rect 35020 47300 35076 47356
rect 35076 47300 35080 47356
rect 35016 47296 35080 47300
rect 35096 47356 35160 47360
rect 35096 47300 35100 47356
rect 35100 47300 35156 47356
rect 35156 47300 35160 47356
rect 35096 47296 35160 47300
rect 35176 47356 35240 47360
rect 35176 47300 35180 47356
rect 35180 47300 35236 47356
rect 35236 47300 35240 47356
rect 35176 47296 35240 47300
rect 19576 46812 19640 46816
rect 19576 46756 19580 46812
rect 19580 46756 19636 46812
rect 19636 46756 19640 46812
rect 19576 46752 19640 46756
rect 19656 46812 19720 46816
rect 19656 46756 19660 46812
rect 19660 46756 19716 46812
rect 19716 46756 19720 46812
rect 19656 46752 19720 46756
rect 19736 46812 19800 46816
rect 19736 46756 19740 46812
rect 19740 46756 19796 46812
rect 19796 46756 19800 46812
rect 19736 46752 19800 46756
rect 19816 46812 19880 46816
rect 19816 46756 19820 46812
rect 19820 46756 19876 46812
rect 19876 46756 19880 46812
rect 19816 46752 19880 46756
rect 50296 46812 50360 46816
rect 50296 46756 50300 46812
rect 50300 46756 50356 46812
rect 50356 46756 50360 46812
rect 50296 46752 50360 46756
rect 50376 46812 50440 46816
rect 50376 46756 50380 46812
rect 50380 46756 50436 46812
rect 50436 46756 50440 46812
rect 50376 46752 50440 46756
rect 50456 46812 50520 46816
rect 50456 46756 50460 46812
rect 50460 46756 50516 46812
rect 50516 46756 50520 46812
rect 50456 46752 50520 46756
rect 50536 46812 50600 46816
rect 50536 46756 50540 46812
rect 50540 46756 50596 46812
rect 50596 46756 50600 46812
rect 50536 46752 50600 46756
rect 4216 46268 4280 46272
rect 4216 46212 4220 46268
rect 4220 46212 4276 46268
rect 4276 46212 4280 46268
rect 4216 46208 4280 46212
rect 4296 46268 4360 46272
rect 4296 46212 4300 46268
rect 4300 46212 4356 46268
rect 4356 46212 4360 46268
rect 4296 46208 4360 46212
rect 4376 46268 4440 46272
rect 4376 46212 4380 46268
rect 4380 46212 4436 46268
rect 4436 46212 4440 46268
rect 4376 46208 4440 46212
rect 4456 46268 4520 46272
rect 4456 46212 4460 46268
rect 4460 46212 4516 46268
rect 4516 46212 4520 46268
rect 4456 46208 4520 46212
rect 34936 46268 35000 46272
rect 34936 46212 34940 46268
rect 34940 46212 34996 46268
rect 34996 46212 35000 46268
rect 34936 46208 35000 46212
rect 35016 46268 35080 46272
rect 35016 46212 35020 46268
rect 35020 46212 35076 46268
rect 35076 46212 35080 46268
rect 35016 46208 35080 46212
rect 35096 46268 35160 46272
rect 35096 46212 35100 46268
rect 35100 46212 35156 46268
rect 35156 46212 35160 46268
rect 35096 46208 35160 46212
rect 35176 46268 35240 46272
rect 35176 46212 35180 46268
rect 35180 46212 35236 46268
rect 35236 46212 35240 46268
rect 35176 46208 35240 46212
rect 19576 45724 19640 45728
rect 19576 45668 19580 45724
rect 19580 45668 19636 45724
rect 19636 45668 19640 45724
rect 19576 45664 19640 45668
rect 19656 45724 19720 45728
rect 19656 45668 19660 45724
rect 19660 45668 19716 45724
rect 19716 45668 19720 45724
rect 19656 45664 19720 45668
rect 19736 45724 19800 45728
rect 19736 45668 19740 45724
rect 19740 45668 19796 45724
rect 19796 45668 19800 45724
rect 19736 45664 19800 45668
rect 19816 45724 19880 45728
rect 19816 45668 19820 45724
rect 19820 45668 19876 45724
rect 19876 45668 19880 45724
rect 19816 45664 19880 45668
rect 50296 45724 50360 45728
rect 50296 45668 50300 45724
rect 50300 45668 50356 45724
rect 50356 45668 50360 45724
rect 50296 45664 50360 45668
rect 50376 45724 50440 45728
rect 50376 45668 50380 45724
rect 50380 45668 50436 45724
rect 50436 45668 50440 45724
rect 50376 45664 50440 45668
rect 50456 45724 50520 45728
rect 50456 45668 50460 45724
rect 50460 45668 50516 45724
rect 50516 45668 50520 45724
rect 50456 45664 50520 45668
rect 50536 45724 50600 45728
rect 50536 45668 50540 45724
rect 50540 45668 50596 45724
rect 50596 45668 50600 45724
rect 50536 45664 50600 45668
rect 4216 45180 4280 45184
rect 4216 45124 4220 45180
rect 4220 45124 4276 45180
rect 4276 45124 4280 45180
rect 4216 45120 4280 45124
rect 4296 45180 4360 45184
rect 4296 45124 4300 45180
rect 4300 45124 4356 45180
rect 4356 45124 4360 45180
rect 4296 45120 4360 45124
rect 4376 45180 4440 45184
rect 4376 45124 4380 45180
rect 4380 45124 4436 45180
rect 4436 45124 4440 45180
rect 4376 45120 4440 45124
rect 4456 45180 4520 45184
rect 4456 45124 4460 45180
rect 4460 45124 4516 45180
rect 4516 45124 4520 45180
rect 4456 45120 4520 45124
rect 34936 45180 35000 45184
rect 34936 45124 34940 45180
rect 34940 45124 34996 45180
rect 34996 45124 35000 45180
rect 34936 45120 35000 45124
rect 35016 45180 35080 45184
rect 35016 45124 35020 45180
rect 35020 45124 35076 45180
rect 35076 45124 35080 45180
rect 35016 45120 35080 45124
rect 35096 45180 35160 45184
rect 35096 45124 35100 45180
rect 35100 45124 35156 45180
rect 35156 45124 35160 45180
rect 35096 45120 35160 45124
rect 35176 45180 35240 45184
rect 35176 45124 35180 45180
rect 35180 45124 35236 45180
rect 35236 45124 35240 45180
rect 35176 45120 35240 45124
rect 19576 44636 19640 44640
rect 19576 44580 19580 44636
rect 19580 44580 19636 44636
rect 19636 44580 19640 44636
rect 19576 44576 19640 44580
rect 19656 44636 19720 44640
rect 19656 44580 19660 44636
rect 19660 44580 19716 44636
rect 19716 44580 19720 44636
rect 19656 44576 19720 44580
rect 19736 44636 19800 44640
rect 19736 44580 19740 44636
rect 19740 44580 19796 44636
rect 19796 44580 19800 44636
rect 19736 44576 19800 44580
rect 19816 44636 19880 44640
rect 19816 44580 19820 44636
rect 19820 44580 19876 44636
rect 19876 44580 19880 44636
rect 19816 44576 19880 44580
rect 50296 44636 50360 44640
rect 50296 44580 50300 44636
rect 50300 44580 50356 44636
rect 50356 44580 50360 44636
rect 50296 44576 50360 44580
rect 50376 44636 50440 44640
rect 50376 44580 50380 44636
rect 50380 44580 50436 44636
rect 50436 44580 50440 44636
rect 50376 44576 50440 44580
rect 50456 44636 50520 44640
rect 50456 44580 50460 44636
rect 50460 44580 50516 44636
rect 50516 44580 50520 44636
rect 50456 44576 50520 44580
rect 50536 44636 50600 44640
rect 50536 44580 50540 44636
rect 50540 44580 50596 44636
rect 50596 44580 50600 44636
rect 50536 44576 50600 44580
rect 4216 44092 4280 44096
rect 4216 44036 4220 44092
rect 4220 44036 4276 44092
rect 4276 44036 4280 44092
rect 4216 44032 4280 44036
rect 4296 44092 4360 44096
rect 4296 44036 4300 44092
rect 4300 44036 4356 44092
rect 4356 44036 4360 44092
rect 4296 44032 4360 44036
rect 4376 44092 4440 44096
rect 4376 44036 4380 44092
rect 4380 44036 4436 44092
rect 4436 44036 4440 44092
rect 4376 44032 4440 44036
rect 4456 44092 4520 44096
rect 4456 44036 4460 44092
rect 4460 44036 4516 44092
rect 4516 44036 4520 44092
rect 4456 44032 4520 44036
rect 34936 44092 35000 44096
rect 34936 44036 34940 44092
rect 34940 44036 34996 44092
rect 34996 44036 35000 44092
rect 34936 44032 35000 44036
rect 35016 44092 35080 44096
rect 35016 44036 35020 44092
rect 35020 44036 35076 44092
rect 35076 44036 35080 44092
rect 35016 44032 35080 44036
rect 35096 44092 35160 44096
rect 35096 44036 35100 44092
rect 35100 44036 35156 44092
rect 35156 44036 35160 44092
rect 35096 44032 35160 44036
rect 35176 44092 35240 44096
rect 35176 44036 35180 44092
rect 35180 44036 35236 44092
rect 35236 44036 35240 44092
rect 35176 44032 35240 44036
rect 19576 43548 19640 43552
rect 19576 43492 19580 43548
rect 19580 43492 19636 43548
rect 19636 43492 19640 43548
rect 19576 43488 19640 43492
rect 19656 43548 19720 43552
rect 19656 43492 19660 43548
rect 19660 43492 19716 43548
rect 19716 43492 19720 43548
rect 19656 43488 19720 43492
rect 19736 43548 19800 43552
rect 19736 43492 19740 43548
rect 19740 43492 19796 43548
rect 19796 43492 19800 43548
rect 19736 43488 19800 43492
rect 19816 43548 19880 43552
rect 19816 43492 19820 43548
rect 19820 43492 19876 43548
rect 19876 43492 19880 43548
rect 19816 43488 19880 43492
rect 50296 43548 50360 43552
rect 50296 43492 50300 43548
rect 50300 43492 50356 43548
rect 50356 43492 50360 43548
rect 50296 43488 50360 43492
rect 50376 43548 50440 43552
rect 50376 43492 50380 43548
rect 50380 43492 50436 43548
rect 50436 43492 50440 43548
rect 50376 43488 50440 43492
rect 50456 43548 50520 43552
rect 50456 43492 50460 43548
rect 50460 43492 50516 43548
rect 50516 43492 50520 43548
rect 50456 43488 50520 43492
rect 50536 43548 50600 43552
rect 50536 43492 50540 43548
rect 50540 43492 50596 43548
rect 50596 43492 50600 43548
rect 50536 43488 50600 43492
rect 4216 43004 4280 43008
rect 4216 42948 4220 43004
rect 4220 42948 4276 43004
rect 4276 42948 4280 43004
rect 4216 42944 4280 42948
rect 4296 43004 4360 43008
rect 4296 42948 4300 43004
rect 4300 42948 4356 43004
rect 4356 42948 4360 43004
rect 4296 42944 4360 42948
rect 4376 43004 4440 43008
rect 4376 42948 4380 43004
rect 4380 42948 4436 43004
rect 4436 42948 4440 43004
rect 4376 42944 4440 42948
rect 4456 43004 4520 43008
rect 4456 42948 4460 43004
rect 4460 42948 4516 43004
rect 4516 42948 4520 43004
rect 4456 42944 4520 42948
rect 34936 43004 35000 43008
rect 34936 42948 34940 43004
rect 34940 42948 34996 43004
rect 34996 42948 35000 43004
rect 34936 42944 35000 42948
rect 35016 43004 35080 43008
rect 35016 42948 35020 43004
rect 35020 42948 35076 43004
rect 35076 42948 35080 43004
rect 35016 42944 35080 42948
rect 35096 43004 35160 43008
rect 35096 42948 35100 43004
rect 35100 42948 35156 43004
rect 35156 42948 35160 43004
rect 35096 42944 35160 42948
rect 35176 43004 35240 43008
rect 35176 42948 35180 43004
rect 35180 42948 35236 43004
rect 35236 42948 35240 43004
rect 35176 42944 35240 42948
rect 19576 42460 19640 42464
rect 19576 42404 19580 42460
rect 19580 42404 19636 42460
rect 19636 42404 19640 42460
rect 19576 42400 19640 42404
rect 19656 42460 19720 42464
rect 19656 42404 19660 42460
rect 19660 42404 19716 42460
rect 19716 42404 19720 42460
rect 19656 42400 19720 42404
rect 19736 42460 19800 42464
rect 19736 42404 19740 42460
rect 19740 42404 19796 42460
rect 19796 42404 19800 42460
rect 19736 42400 19800 42404
rect 19816 42460 19880 42464
rect 19816 42404 19820 42460
rect 19820 42404 19876 42460
rect 19876 42404 19880 42460
rect 19816 42400 19880 42404
rect 50296 42460 50360 42464
rect 50296 42404 50300 42460
rect 50300 42404 50356 42460
rect 50356 42404 50360 42460
rect 50296 42400 50360 42404
rect 50376 42460 50440 42464
rect 50376 42404 50380 42460
rect 50380 42404 50436 42460
rect 50436 42404 50440 42460
rect 50376 42400 50440 42404
rect 50456 42460 50520 42464
rect 50456 42404 50460 42460
rect 50460 42404 50516 42460
rect 50516 42404 50520 42460
rect 50456 42400 50520 42404
rect 50536 42460 50600 42464
rect 50536 42404 50540 42460
rect 50540 42404 50596 42460
rect 50596 42404 50600 42460
rect 50536 42400 50600 42404
rect 4216 41916 4280 41920
rect 4216 41860 4220 41916
rect 4220 41860 4276 41916
rect 4276 41860 4280 41916
rect 4216 41856 4280 41860
rect 4296 41916 4360 41920
rect 4296 41860 4300 41916
rect 4300 41860 4356 41916
rect 4356 41860 4360 41916
rect 4296 41856 4360 41860
rect 4376 41916 4440 41920
rect 4376 41860 4380 41916
rect 4380 41860 4436 41916
rect 4436 41860 4440 41916
rect 4376 41856 4440 41860
rect 4456 41916 4520 41920
rect 4456 41860 4460 41916
rect 4460 41860 4516 41916
rect 4516 41860 4520 41916
rect 4456 41856 4520 41860
rect 34936 41916 35000 41920
rect 34936 41860 34940 41916
rect 34940 41860 34996 41916
rect 34996 41860 35000 41916
rect 34936 41856 35000 41860
rect 35016 41916 35080 41920
rect 35016 41860 35020 41916
rect 35020 41860 35076 41916
rect 35076 41860 35080 41916
rect 35016 41856 35080 41860
rect 35096 41916 35160 41920
rect 35096 41860 35100 41916
rect 35100 41860 35156 41916
rect 35156 41860 35160 41916
rect 35096 41856 35160 41860
rect 35176 41916 35240 41920
rect 35176 41860 35180 41916
rect 35180 41860 35236 41916
rect 35236 41860 35240 41916
rect 35176 41856 35240 41860
rect 19576 41372 19640 41376
rect 19576 41316 19580 41372
rect 19580 41316 19636 41372
rect 19636 41316 19640 41372
rect 19576 41312 19640 41316
rect 19656 41372 19720 41376
rect 19656 41316 19660 41372
rect 19660 41316 19716 41372
rect 19716 41316 19720 41372
rect 19656 41312 19720 41316
rect 19736 41372 19800 41376
rect 19736 41316 19740 41372
rect 19740 41316 19796 41372
rect 19796 41316 19800 41372
rect 19736 41312 19800 41316
rect 19816 41372 19880 41376
rect 19816 41316 19820 41372
rect 19820 41316 19876 41372
rect 19876 41316 19880 41372
rect 19816 41312 19880 41316
rect 50296 41372 50360 41376
rect 50296 41316 50300 41372
rect 50300 41316 50356 41372
rect 50356 41316 50360 41372
rect 50296 41312 50360 41316
rect 50376 41372 50440 41376
rect 50376 41316 50380 41372
rect 50380 41316 50436 41372
rect 50436 41316 50440 41372
rect 50376 41312 50440 41316
rect 50456 41372 50520 41376
rect 50456 41316 50460 41372
rect 50460 41316 50516 41372
rect 50516 41316 50520 41372
rect 50456 41312 50520 41316
rect 50536 41372 50600 41376
rect 50536 41316 50540 41372
rect 50540 41316 50596 41372
rect 50596 41316 50600 41372
rect 50536 41312 50600 41316
rect 4216 40828 4280 40832
rect 4216 40772 4220 40828
rect 4220 40772 4276 40828
rect 4276 40772 4280 40828
rect 4216 40768 4280 40772
rect 4296 40828 4360 40832
rect 4296 40772 4300 40828
rect 4300 40772 4356 40828
rect 4356 40772 4360 40828
rect 4296 40768 4360 40772
rect 4376 40828 4440 40832
rect 4376 40772 4380 40828
rect 4380 40772 4436 40828
rect 4436 40772 4440 40828
rect 4376 40768 4440 40772
rect 4456 40828 4520 40832
rect 4456 40772 4460 40828
rect 4460 40772 4516 40828
rect 4516 40772 4520 40828
rect 4456 40768 4520 40772
rect 34936 40828 35000 40832
rect 34936 40772 34940 40828
rect 34940 40772 34996 40828
rect 34996 40772 35000 40828
rect 34936 40768 35000 40772
rect 35016 40828 35080 40832
rect 35016 40772 35020 40828
rect 35020 40772 35076 40828
rect 35076 40772 35080 40828
rect 35016 40768 35080 40772
rect 35096 40828 35160 40832
rect 35096 40772 35100 40828
rect 35100 40772 35156 40828
rect 35156 40772 35160 40828
rect 35096 40768 35160 40772
rect 35176 40828 35240 40832
rect 35176 40772 35180 40828
rect 35180 40772 35236 40828
rect 35236 40772 35240 40828
rect 35176 40768 35240 40772
rect 19576 40284 19640 40288
rect 19576 40228 19580 40284
rect 19580 40228 19636 40284
rect 19636 40228 19640 40284
rect 19576 40224 19640 40228
rect 19656 40284 19720 40288
rect 19656 40228 19660 40284
rect 19660 40228 19716 40284
rect 19716 40228 19720 40284
rect 19656 40224 19720 40228
rect 19736 40284 19800 40288
rect 19736 40228 19740 40284
rect 19740 40228 19796 40284
rect 19796 40228 19800 40284
rect 19736 40224 19800 40228
rect 19816 40284 19880 40288
rect 19816 40228 19820 40284
rect 19820 40228 19876 40284
rect 19876 40228 19880 40284
rect 19816 40224 19880 40228
rect 50296 40284 50360 40288
rect 50296 40228 50300 40284
rect 50300 40228 50356 40284
rect 50356 40228 50360 40284
rect 50296 40224 50360 40228
rect 50376 40284 50440 40288
rect 50376 40228 50380 40284
rect 50380 40228 50436 40284
rect 50436 40228 50440 40284
rect 50376 40224 50440 40228
rect 50456 40284 50520 40288
rect 50456 40228 50460 40284
rect 50460 40228 50516 40284
rect 50516 40228 50520 40284
rect 50456 40224 50520 40228
rect 50536 40284 50600 40288
rect 50536 40228 50540 40284
rect 50540 40228 50596 40284
rect 50596 40228 50600 40284
rect 50536 40224 50600 40228
rect 4216 39740 4280 39744
rect 4216 39684 4220 39740
rect 4220 39684 4276 39740
rect 4276 39684 4280 39740
rect 4216 39680 4280 39684
rect 4296 39740 4360 39744
rect 4296 39684 4300 39740
rect 4300 39684 4356 39740
rect 4356 39684 4360 39740
rect 4296 39680 4360 39684
rect 4376 39740 4440 39744
rect 4376 39684 4380 39740
rect 4380 39684 4436 39740
rect 4436 39684 4440 39740
rect 4376 39680 4440 39684
rect 4456 39740 4520 39744
rect 4456 39684 4460 39740
rect 4460 39684 4516 39740
rect 4516 39684 4520 39740
rect 4456 39680 4520 39684
rect 34936 39740 35000 39744
rect 34936 39684 34940 39740
rect 34940 39684 34996 39740
rect 34996 39684 35000 39740
rect 34936 39680 35000 39684
rect 35016 39740 35080 39744
rect 35016 39684 35020 39740
rect 35020 39684 35076 39740
rect 35076 39684 35080 39740
rect 35016 39680 35080 39684
rect 35096 39740 35160 39744
rect 35096 39684 35100 39740
rect 35100 39684 35156 39740
rect 35156 39684 35160 39740
rect 35096 39680 35160 39684
rect 35176 39740 35240 39744
rect 35176 39684 35180 39740
rect 35180 39684 35236 39740
rect 35236 39684 35240 39740
rect 35176 39680 35240 39684
rect 19576 39196 19640 39200
rect 19576 39140 19580 39196
rect 19580 39140 19636 39196
rect 19636 39140 19640 39196
rect 19576 39136 19640 39140
rect 19656 39196 19720 39200
rect 19656 39140 19660 39196
rect 19660 39140 19716 39196
rect 19716 39140 19720 39196
rect 19656 39136 19720 39140
rect 19736 39196 19800 39200
rect 19736 39140 19740 39196
rect 19740 39140 19796 39196
rect 19796 39140 19800 39196
rect 19736 39136 19800 39140
rect 19816 39196 19880 39200
rect 19816 39140 19820 39196
rect 19820 39140 19876 39196
rect 19876 39140 19880 39196
rect 19816 39136 19880 39140
rect 50296 39196 50360 39200
rect 50296 39140 50300 39196
rect 50300 39140 50356 39196
rect 50356 39140 50360 39196
rect 50296 39136 50360 39140
rect 50376 39196 50440 39200
rect 50376 39140 50380 39196
rect 50380 39140 50436 39196
rect 50436 39140 50440 39196
rect 50376 39136 50440 39140
rect 50456 39196 50520 39200
rect 50456 39140 50460 39196
rect 50460 39140 50516 39196
rect 50516 39140 50520 39196
rect 50456 39136 50520 39140
rect 50536 39196 50600 39200
rect 50536 39140 50540 39196
rect 50540 39140 50596 39196
rect 50596 39140 50600 39196
rect 50536 39136 50600 39140
rect 4216 38652 4280 38656
rect 4216 38596 4220 38652
rect 4220 38596 4276 38652
rect 4276 38596 4280 38652
rect 4216 38592 4280 38596
rect 4296 38652 4360 38656
rect 4296 38596 4300 38652
rect 4300 38596 4356 38652
rect 4356 38596 4360 38652
rect 4296 38592 4360 38596
rect 4376 38652 4440 38656
rect 4376 38596 4380 38652
rect 4380 38596 4436 38652
rect 4436 38596 4440 38652
rect 4376 38592 4440 38596
rect 4456 38652 4520 38656
rect 4456 38596 4460 38652
rect 4460 38596 4516 38652
rect 4516 38596 4520 38652
rect 4456 38592 4520 38596
rect 34936 38652 35000 38656
rect 34936 38596 34940 38652
rect 34940 38596 34996 38652
rect 34996 38596 35000 38652
rect 34936 38592 35000 38596
rect 35016 38652 35080 38656
rect 35016 38596 35020 38652
rect 35020 38596 35076 38652
rect 35076 38596 35080 38652
rect 35016 38592 35080 38596
rect 35096 38652 35160 38656
rect 35096 38596 35100 38652
rect 35100 38596 35156 38652
rect 35156 38596 35160 38652
rect 35096 38592 35160 38596
rect 35176 38652 35240 38656
rect 35176 38596 35180 38652
rect 35180 38596 35236 38652
rect 35236 38596 35240 38652
rect 35176 38592 35240 38596
rect 19576 38108 19640 38112
rect 19576 38052 19580 38108
rect 19580 38052 19636 38108
rect 19636 38052 19640 38108
rect 19576 38048 19640 38052
rect 19656 38108 19720 38112
rect 19656 38052 19660 38108
rect 19660 38052 19716 38108
rect 19716 38052 19720 38108
rect 19656 38048 19720 38052
rect 19736 38108 19800 38112
rect 19736 38052 19740 38108
rect 19740 38052 19796 38108
rect 19796 38052 19800 38108
rect 19736 38048 19800 38052
rect 19816 38108 19880 38112
rect 19816 38052 19820 38108
rect 19820 38052 19876 38108
rect 19876 38052 19880 38108
rect 19816 38048 19880 38052
rect 50296 38108 50360 38112
rect 50296 38052 50300 38108
rect 50300 38052 50356 38108
rect 50356 38052 50360 38108
rect 50296 38048 50360 38052
rect 50376 38108 50440 38112
rect 50376 38052 50380 38108
rect 50380 38052 50436 38108
rect 50436 38052 50440 38108
rect 50376 38048 50440 38052
rect 50456 38108 50520 38112
rect 50456 38052 50460 38108
rect 50460 38052 50516 38108
rect 50516 38052 50520 38108
rect 50456 38048 50520 38052
rect 50536 38108 50600 38112
rect 50536 38052 50540 38108
rect 50540 38052 50596 38108
rect 50596 38052 50600 38108
rect 50536 38048 50600 38052
rect 4216 37564 4280 37568
rect 4216 37508 4220 37564
rect 4220 37508 4276 37564
rect 4276 37508 4280 37564
rect 4216 37504 4280 37508
rect 4296 37564 4360 37568
rect 4296 37508 4300 37564
rect 4300 37508 4356 37564
rect 4356 37508 4360 37564
rect 4296 37504 4360 37508
rect 4376 37564 4440 37568
rect 4376 37508 4380 37564
rect 4380 37508 4436 37564
rect 4436 37508 4440 37564
rect 4376 37504 4440 37508
rect 4456 37564 4520 37568
rect 4456 37508 4460 37564
rect 4460 37508 4516 37564
rect 4516 37508 4520 37564
rect 4456 37504 4520 37508
rect 34936 37564 35000 37568
rect 34936 37508 34940 37564
rect 34940 37508 34996 37564
rect 34996 37508 35000 37564
rect 34936 37504 35000 37508
rect 35016 37564 35080 37568
rect 35016 37508 35020 37564
rect 35020 37508 35076 37564
rect 35076 37508 35080 37564
rect 35016 37504 35080 37508
rect 35096 37564 35160 37568
rect 35096 37508 35100 37564
rect 35100 37508 35156 37564
rect 35156 37508 35160 37564
rect 35096 37504 35160 37508
rect 35176 37564 35240 37568
rect 35176 37508 35180 37564
rect 35180 37508 35236 37564
rect 35236 37508 35240 37564
rect 35176 37504 35240 37508
rect 19576 37020 19640 37024
rect 19576 36964 19580 37020
rect 19580 36964 19636 37020
rect 19636 36964 19640 37020
rect 19576 36960 19640 36964
rect 19656 37020 19720 37024
rect 19656 36964 19660 37020
rect 19660 36964 19716 37020
rect 19716 36964 19720 37020
rect 19656 36960 19720 36964
rect 19736 37020 19800 37024
rect 19736 36964 19740 37020
rect 19740 36964 19796 37020
rect 19796 36964 19800 37020
rect 19736 36960 19800 36964
rect 19816 37020 19880 37024
rect 19816 36964 19820 37020
rect 19820 36964 19876 37020
rect 19876 36964 19880 37020
rect 19816 36960 19880 36964
rect 50296 37020 50360 37024
rect 50296 36964 50300 37020
rect 50300 36964 50356 37020
rect 50356 36964 50360 37020
rect 50296 36960 50360 36964
rect 50376 37020 50440 37024
rect 50376 36964 50380 37020
rect 50380 36964 50436 37020
rect 50436 36964 50440 37020
rect 50376 36960 50440 36964
rect 50456 37020 50520 37024
rect 50456 36964 50460 37020
rect 50460 36964 50516 37020
rect 50516 36964 50520 37020
rect 50456 36960 50520 36964
rect 50536 37020 50600 37024
rect 50536 36964 50540 37020
rect 50540 36964 50596 37020
rect 50596 36964 50600 37020
rect 50536 36960 50600 36964
rect 4216 36476 4280 36480
rect 4216 36420 4220 36476
rect 4220 36420 4276 36476
rect 4276 36420 4280 36476
rect 4216 36416 4280 36420
rect 4296 36476 4360 36480
rect 4296 36420 4300 36476
rect 4300 36420 4356 36476
rect 4356 36420 4360 36476
rect 4296 36416 4360 36420
rect 4376 36476 4440 36480
rect 4376 36420 4380 36476
rect 4380 36420 4436 36476
rect 4436 36420 4440 36476
rect 4376 36416 4440 36420
rect 4456 36476 4520 36480
rect 4456 36420 4460 36476
rect 4460 36420 4516 36476
rect 4516 36420 4520 36476
rect 4456 36416 4520 36420
rect 34936 36476 35000 36480
rect 34936 36420 34940 36476
rect 34940 36420 34996 36476
rect 34996 36420 35000 36476
rect 34936 36416 35000 36420
rect 35016 36476 35080 36480
rect 35016 36420 35020 36476
rect 35020 36420 35076 36476
rect 35076 36420 35080 36476
rect 35016 36416 35080 36420
rect 35096 36476 35160 36480
rect 35096 36420 35100 36476
rect 35100 36420 35156 36476
rect 35156 36420 35160 36476
rect 35096 36416 35160 36420
rect 35176 36476 35240 36480
rect 35176 36420 35180 36476
rect 35180 36420 35236 36476
rect 35236 36420 35240 36476
rect 35176 36416 35240 36420
rect 19576 35932 19640 35936
rect 19576 35876 19580 35932
rect 19580 35876 19636 35932
rect 19636 35876 19640 35932
rect 19576 35872 19640 35876
rect 19656 35932 19720 35936
rect 19656 35876 19660 35932
rect 19660 35876 19716 35932
rect 19716 35876 19720 35932
rect 19656 35872 19720 35876
rect 19736 35932 19800 35936
rect 19736 35876 19740 35932
rect 19740 35876 19796 35932
rect 19796 35876 19800 35932
rect 19736 35872 19800 35876
rect 19816 35932 19880 35936
rect 19816 35876 19820 35932
rect 19820 35876 19876 35932
rect 19876 35876 19880 35932
rect 19816 35872 19880 35876
rect 50296 35932 50360 35936
rect 50296 35876 50300 35932
rect 50300 35876 50356 35932
rect 50356 35876 50360 35932
rect 50296 35872 50360 35876
rect 50376 35932 50440 35936
rect 50376 35876 50380 35932
rect 50380 35876 50436 35932
rect 50436 35876 50440 35932
rect 50376 35872 50440 35876
rect 50456 35932 50520 35936
rect 50456 35876 50460 35932
rect 50460 35876 50516 35932
rect 50516 35876 50520 35932
rect 50456 35872 50520 35876
rect 50536 35932 50600 35936
rect 50536 35876 50540 35932
rect 50540 35876 50596 35932
rect 50596 35876 50600 35932
rect 50536 35872 50600 35876
rect 4216 35388 4280 35392
rect 4216 35332 4220 35388
rect 4220 35332 4276 35388
rect 4276 35332 4280 35388
rect 4216 35328 4280 35332
rect 4296 35388 4360 35392
rect 4296 35332 4300 35388
rect 4300 35332 4356 35388
rect 4356 35332 4360 35388
rect 4296 35328 4360 35332
rect 4376 35388 4440 35392
rect 4376 35332 4380 35388
rect 4380 35332 4436 35388
rect 4436 35332 4440 35388
rect 4376 35328 4440 35332
rect 4456 35388 4520 35392
rect 4456 35332 4460 35388
rect 4460 35332 4516 35388
rect 4516 35332 4520 35388
rect 4456 35328 4520 35332
rect 34936 35388 35000 35392
rect 34936 35332 34940 35388
rect 34940 35332 34996 35388
rect 34996 35332 35000 35388
rect 34936 35328 35000 35332
rect 35016 35388 35080 35392
rect 35016 35332 35020 35388
rect 35020 35332 35076 35388
rect 35076 35332 35080 35388
rect 35016 35328 35080 35332
rect 35096 35388 35160 35392
rect 35096 35332 35100 35388
rect 35100 35332 35156 35388
rect 35156 35332 35160 35388
rect 35096 35328 35160 35332
rect 35176 35388 35240 35392
rect 35176 35332 35180 35388
rect 35180 35332 35236 35388
rect 35236 35332 35240 35388
rect 35176 35328 35240 35332
rect 19576 34844 19640 34848
rect 19576 34788 19580 34844
rect 19580 34788 19636 34844
rect 19636 34788 19640 34844
rect 19576 34784 19640 34788
rect 19656 34844 19720 34848
rect 19656 34788 19660 34844
rect 19660 34788 19716 34844
rect 19716 34788 19720 34844
rect 19656 34784 19720 34788
rect 19736 34844 19800 34848
rect 19736 34788 19740 34844
rect 19740 34788 19796 34844
rect 19796 34788 19800 34844
rect 19736 34784 19800 34788
rect 19816 34844 19880 34848
rect 19816 34788 19820 34844
rect 19820 34788 19876 34844
rect 19876 34788 19880 34844
rect 19816 34784 19880 34788
rect 50296 34844 50360 34848
rect 50296 34788 50300 34844
rect 50300 34788 50356 34844
rect 50356 34788 50360 34844
rect 50296 34784 50360 34788
rect 50376 34844 50440 34848
rect 50376 34788 50380 34844
rect 50380 34788 50436 34844
rect 50436 34788 50440 34844
rect 50376 34784 50440 34788
rect 50456 34844 50520 34848
rect 50456 34788 50460 34844
rect 50460 34788 50516 34844
rect 50516 34788 50520 34844
rect 50456 34784 50520 34788
rect 50536 34844 50600 34848
rect 50536 34788 50540 34844
rect 50540 34788 50596 34844
rect 50596 34788 50600 34844
rect 50536 34784 50600 34788
rect 4216 34300 4280 34304
rect 4216 34244 4220 34300
rect 4220 34244 4276 34300
rect 4276 34244 4280 34300
rect 4216 34240 4280 34244
rect 4296 34300 4360 34304
rect 4296 34244 4300 34300
rect 4300 34244 4356 34300
rect 4356 34244 4360 34300
rect 4296 34240 4360 34244
rect 4376 34300 4440 34304
rect 4376 34244 4380 34300
rect 4380 34244 4436 34300
rect 4436 34244 4440 34300
rect 4376 34240 4440 34244
rect 4456 34300 4520 34304
rect 4456 34244 4460 34300
rect 4460 34244 4516 34300
rect 4516 34244 4520 34300
rect 4456 34240 4520 34244
rect 34936 34300 35000 34304
rect 34936 34244 34940 34300
rect 34940 34244 34996 34300
rect 34996 34244 35000 34300
rect 34936 34240 35000 34244
rect 35016 34300 35080 34304
rect 35016 34244 35020 34300
rect 35020 34244 35076 34300
rect 35076 34244 35080 34300
rect 35016 34240 35080 34244
rect 35096 34300 35160 34304
rect 35096 34244 35100 34300
rect 35100 34244 35156 34300
rect 35156 34244 35160 34300
rect 35096 34240 35160 34244
rect 35176 34300 35240 34304
rect 35176 34244 35180 34300
rect 35180 34244 35236 34300
rect 35236 34244 35240 34300
rect 35176 34240 35240 34244
rect 19576 33756 19640 33760
rect 19576 33700 19580 33756
rect 19580 33700 19636 33756
rect 19636 33700 19640 33756
rect 19576 33696 19640 33700
rect 19656 33756 19720 33760
rect 19656 33700 19660 33756
rect 19660 33700 19716 33756
rect 19716 33700 19720 33756
rect 19656 33696 19720 33700
rect 19736 33756 19800 33760
rect 19736 33700 19740 33756
rect 19740 33700 19796 33756
rect 19796 33700 19800 33756
rect 19736 33696 19800 33700
rect 19816 33756 19880 33760
rect 19816 33700 19820 33756
rect 19820 33700 19876 33756
rect 19876 33700 19880 33756
rect 19816 33696 19880 33700
rect 50296 33756 50360 33760
rect 50296 33700 50300 33756
rect 50300 33700 50356 33756
rect 50356 33700 50360 33756
rect 50296 33696 50360 33700
rect 50376 33756 50440 33760
rect 50376 33700 50380 33756
rect 50380 33700 50436 33756
rect 50436 33700 50440 33756
rect 50376 33696 50440 33700
rect 50456 33756 50520 33760
rect 50456 33700 50460 33756
rect 50460 33700 50516 33756
rect 50516 33700 50520 33756
rect 50456 33696 50520 33700
rect 50536 33756 50600 33760
rect 50536 33700 50540 33756
rect 50540 33700 50596 33756
rect 50596 33700 50600 33756
rect 50536 33696 50600 33700
rect 4216 33212 4280 33216
rect 4216 33156 4220 33212
rect 4220 33156 4276 33212
rect 4276 33156 4280 33212
rect 4216 33152 4280 33156
rect 4296 33212 4360 33216
rect 4296 33156 4300 33212
rect 4300 33156 4356 33212
rect 4356 33156 4360 33212
rect 4296 33152 4360 33156
rect 4376 33212 4440 33216
rect 4376 33156 4380 33212
rect 4380 33156 4436 33212
rect 4436 33156 4440 33212
rect 4376 33152 4440 33156
rect 4456 33212 4520 33216
rect 4456 33156 4460 33212
rect 4460 33156 4516 33212
rect 4516 33156 4520 33212
rect 4456 33152 4520 33156
rect 34936 33212 35000 33216
rect 34936 33156 34940 33212
rect 34940 33156 34996 33212
rect 34996 33156 35000 33212
rect 34936 33152 35000 33156
rect 35016 33212 35080 33216
rect 35016 33156 35020 33212
rect 35020 33156 35076 33212
rect 35076 33156 35080 33212
rect 35016 33152 35080 33156
rect 35096 33212 35160 33216
rect 35096 33156 35100 33212
rect 35100 33156 35156 33212
rect 35156 33156 35160 33212
rect 35096 33152 35160 33156
rect 35176 33212 35240 33216
rect 35176 33156 35180 33212
rect 35180 33156 35236 33212
rect 35236 33156 35240 33212
rect 35176 33152 35240 33156
rect 19576 32668 19640 32672
rect 19576 32612 19580 32668
rect 19580 32612 19636 32668
rect 19636 32612 19640 32668
rect 19576 32608 19640 32612
rect 19656 32668 19720 32672
rect 19656 32612 19660 32668
rect 19660 32612 19716 32668
rect 19716 32612 19720 32668
rect 19656 32608 19720 32612
rect 19736 32668 19800 32672
rect 19736 32612 19740 32668
rect 19740 32612 19796 32668
rect 19796 32612 19800 32668
rect 19736 32608 19800 32612
rect 19816 32668 19880 32672
rect 19816 32612 19820 32668
rect 19820 32612 19876 32668
rect 19876 32612 19880 32668
rect 19816 32608 19880 32612
rect 50296 32668 50360 32672
rect 50296 32612 50300 32668
rect 50300 32612 50356 32668
rect 50356 32612 50360 32668
rect 50296 32608 50360 32612
rect 50376 32668 50440 32672
rect 50376 32612 50380 32668
rect 50380 32612 50436 32668
rect 50436 32612 50440 32668
rect 50376 32608 50440 32612
rect 50456 32668 50520 32672
rect 50456 32612 50460 32668
rect 50460 32612 50516 32668
rect 50516 32612 50520 32668
rect 50456 32608 50520 32612
rect 50536 32668 50600 32672
rect 50536 32612 50540 32668
rect 50540 32612 50596 32668
rect 50596 32612 50600 32668
rect 50536 32608 50600 32612
rect 4216 32124 4280 32128
rect 4216 32068 4220 32124
rect 4220 32068 4276 32124
rect 4276 32068 4280 32124
rect 4216 32064 4280 32068
rect 4296 32124 4360 32128
rect 4296 32068 4300 32124
rect 4300 32068 4356 32124
rect 4356 32068 4360 32124
rect 4296 32064 4360 32068
rect 4376 32124 4440 32128
rect 4376 32068 4380 32124
rect 4380 32068 4436 32124
rect 4436 32068 4440 32124
rect 4376 32064 4440 32068
rect 4456 32124 4520 32128
rect 4456 32068 4460 32124
rect 4460 32068 4516 32124
rect 4516 32068 4520 32124
rect 4456 32064 4520 32068
rect 34936 32124 35000 32128
rect 34936 32068 34940 32124
rect 34940 32068 34996 32124
rect 34996 32068 35000 32124
rect 34936 32064 35000 32068
rect 35016 32124 35080 32128
rect 35016 32068 35020 32124
rect 35020 32068 35076 32124
rect 35076 32068 35080 32124
rect 35016 32064 35080 32068
rect 35096 32124 35160 32128
rect 35096 32068 35100 32124
rect 35100 32068 35156 32124
rect 35156 32068 35160 32124
rect 35096 32064 35160 32068
rect 35176 32124 35240 32128
rect 35176 32068 35180 32124
rect 35180 32068 35236 32124
rect 35236 32068 35240 32124
rect 35176 32064 35240 32068
rect 19576 31580 19640 31584
rect 19576 31524 19580 31580
rect 19580 31524 19636 31580
rect 19636 31524 19640 31580
rect 19576 31520 19640 31524
rect 19656 31580 19720 31584
rect 19656 31524 19660 31580
rect 19660 31524 19716 31580
rect 19716 31524 19720 31580
rect 19656 31520 19720 31524
rect 19736 31580 19800 31584
rect 19736 31524 19740 31580
rect 19740 31524 19796 31580
rect 19796 31524 19800 31580
rect 19736 31520 19800 31524
rect 19816 31580 19880 31584
rect 19816 31524 19820 31580
rect 19820 31524 19876 31580
rect 19876 31524 19880 31580
rect 19816 31520 19880 31524
rect 50296 31580 50360 31584
rect 50296 31524 50300 31580
rect 50300 31524 50356 31580
rect 50356 31524 50360 31580
rect 50296 31520 50360 31524
rect 50376 31580 50440 31584
rect 50376 31524 50380 31580
rect 50380 31524 50436 31580
rect 50436 31524 50440 31580
rect 50376 31520 50440 31524
rect 50456 31580 50520 31584
rect 50456 31524 50460 31580
rect 50460 31524 50516 31580
rect 50516 31524 50520 31580
rect 50456 31520 50520 31524
rect 50536 31580 50600 31584
rect 50536 31524 50540 31580
rect 50540 31524 50596 31580
rect 50596 31524 50600 31580
rect 50536 31520 50600 31524
rect 4216 31036 4280 31040
rect 4216 30980 4220 31036
rect 4220 30980 4276 31036
rect 4276 30980 4280 31036
rect 4216 30976 4280 30980
rect 4296 31036 4360 31040
rect 4296 30980 4300 31036
rect 4300 30980 4356 31036
rect 4356 30980 4360 31036
rect 4296 30976 4360 30980
rect 4376 31036 4440 31040
rect 4376 30980 4380 31036
rect 4380 30980 4436 31036
rect 4436 30980 4440 31036
rect 4376 30976 4440 30980
rect 4456 31036 4520 31040
rect 4456 30980 4460 31036
rect 4460 30980 4516 31036
rect 4516 30980 4520 31036
rect 4456 30976 4520 30980
rect 34936 31036 35000 31040
rect 34936 30980 34940 31036
rect 34940 30980 34996 31036
rect 34996 30980 35000 31036
rect 34936 30976 35000 30980
rect 35016 31036 35080 31040
rect 35016 30980 35020 31036
rect 35020 30980 35076 31036
rect 35076 30980 35080 31036
rect 35016 30976 35080 30980
rect 35096 31036 35160 31040
rect 35096 30980 35100 31036
rect 35100 30980 35156 31036
rect 35156 30980 35160 31036
rect 35096 30976 35160 30980
rect 35176 31036 35240 31040
rect 35176 30980 35180 31036
rect 35180 30980 35236 31036
rect 35236 30980 35240 31036
rect 35176 30976 35240 30980
rect 19576 30492 19640 30496
rect 19576 30436 19580 30492
rect 19580 30436 19636 30492
rect 19636 30436 19640 30492
rect 19576 30432 19640 30436
rect 19656 30492 19720 30496
rect 19656 30436 19660 30492
rect 19660 30436 19716 30492
rect 19716 30436 19720 30492
rect 19656 30432 19720 30436
rect 19736 30492 19800 30496
rect 19736 30436 19740 30492
rect 19740 30436 19796 30492
rect 19796 30436 19800 30492
rect 19736 30432 19800 30436
rect 19816 30492 19880 30496
rect 19816 30436 19820 30492
rect 19820 30436 19876 30492
rect 19876 30436 19880 30492
rect 19816 30432 19880 30436
rect 50296 30492 50360 30496
rect 50296 30436 50300 30492
rect 50300 30436 50356 30492
rect 50356 30436 50360 30492
rect 50296 30432 50360 30436
rect 50376 30492 50440 30496
rect 50376 30436 50380 30492
rect 50380 30436 50436 30492
rect 50436 30436 50440 30492
rect 50376 30432 50440 30436
rect 50456 30492 50520 30496
rect 50456 30436 50460 30492
rect 50460 30436 50516 30492
rect 50516 30436 50520 30492
rect 50456 30432 50520 30436
rect 50536 30492 50600 30496
rect 50536 30436 50540 30492
rect 50540 30436 50596 30492
rect 50596 30436 50600 30492
rect 50536 30432 50600 30436
rect 4216 29948 4280 29952
rect 4216 29892 4220 29948
rect 4220 29892 4276 29948
rect 4276 29892 4280 29948
rect 4216 29888 4280 29892
rect 4296 29948 4360 29952
rect 4296 29892 4300 29948
rect 4300 29892 4356 29948
rect 4356 29892 4360 29948
rect 4296 29888 4360 29892
rect 4376 29948 4440 29952
rect 4376 29892 4380 29948
rect 4380 29892 4436 29948
rect 4436 29892 4440 29948
rect 4376 29888 4440 29892
rect 4456 29948 4520 29952
rect 4456 29892 4460 29948
rect 4460 29892 4516 29948
rect 4516 29892 4520 29948
rect 4456 29888 4520 29892
rect 34936 29948 35000 29952
rect 34936 29892 34940 29948
rect 34940 29892 34996 29948
rect 34996 29892 35000 29948
rect 34936 29888 35000 29892
rect 35016 29948 35080 29952
rect 35016 29892 35020 29948
rect 35020 29892 35076 29948
rect 35076 29892 35080 29948
rect 35016 29888 35080 29892
rect 35096 29948 35160 29952
rect 35096 29892 35100 29948
rect 35100 29892 35156 29948
rect 35156 29892 35160 29948
rect 35096 29888 35160 29892
rect 35176 29948 35240 29952
rect 35176 29892 35180 29948
rect 35180 29892 35236 29948
rect 35236 29892 35240 29948
rect 35176 29888 35240 29892
rect 19576 29404 19640 29408
rect 19576 29348 19580 29404
rect 19580 29348 19636 29404
rect 19636 29348 19640 29404
rect 19576 29344 19640 29348
rect 19656 29404 19720 29408
rect 19656 29348 19660 29404
rect 19660 29348 19716 29404
rect 19716 29348 19720 29404
rect 19656 29344 19720 29348
rect 19736 29404 19800 29408
rect 19736 29348 19740 29404
rect 19740 29348 19796 29404
rect 19796 29348 19800 29404
rect 19736 29344 19800 29348
rect 19816 29404 19880 29408
rect 19816 29348 19820 29404
rect 19820 29348 19876 29404
rect 19876 29348 19880 29404
rect 19816 29344 19880 29348
rect 50296 29404 50360 29408
rect 50296 29348 50300 29404
rect 50300 29348 50356 29404
rect 50356 29348 50360 29404
rect 50296 29344 50360 29348
rect 50376 29404 50440 29408
rect 50376 29348 50380 29404
rect 50380 29348 50436 29404
rect 50436 29348 50440 29404
rect 50376 29344 50440 29348
rect 50456 29404 50520 29408
rect 50456 29348 50460 29404
rect 50460 29348 50516 29404
rect 50516 29348 50520 29404
rect 50456 29344 50520 29348
rect 50536 29404 50600 29408
rect 50536 29348 50540 29404
rect 50540 29348 50596 29404
rect 50596 29348 50600 29404
rect 50536 29344 50600 29348
rect 4216 28860 4280 28864
rect 4216 28804 4220 28860
rect 4220 28804 4276 28860
rect 4276 28804 4280 28860
rect 4216 28800 4280 28804
rect 4296 28860 4360 28864
rect 4296 28804 4300 28860
rect 4300 28804 4356 28860
rect 4356 28804 4360 28860
rect 4296 28800 4360 28804
rect 4376 28860 4440 28864
rect 4376 28804 4380 28860
rect 4380 28804 4436 28860
rect 4436 28804 4440 28860
rect 4376 28800 4440 28804
rect 4456 28860 4520 28864
rect 4456 28804 4460 28860
rect 4460 28804 4516 28860
rect 4516 28804 4520 28860
rect 4456 28800 4520 28804
rect 34936 28860 35000 28864
rect 34936 28804 34940 28860
rect 34940 28804 34996 28860
rect 34996 28804 35000 28860
rect 34936 28800 35000 28804
rect 35016 28860 35080 28864
rect 35016 28804 35020 28860
rect 35020 28804 35076 28860
rect 35076 28804 35080 28860
rect 35016 28800 35080 28804
rect 35096 28860 35160 28864
rect 35096 28804 35100 28860
rect 35100 28804 35156 28860
rect 35156 28804 35160 28860
rect 35096 28800 35160 28804
rect 35176 28860 35240 28864
rect 35176 28804 35180 28860
rect 35180 28804 35236 28860
rect 35236 28804 35240 28860
rect 35176 28800 35240 28804
rect 19576 28316 19640 28320
rect 19576 28260 19580 28316
rect 19580 28260 19636 28316
rect 19636 28260 19640 28316
rect 19576 28256 19640 28260
rect 19656 28316 19720 28320
rect 19656 28260 19660 28316
rect 19660 28260 19716 28316
rect 19716 28260 19720 28316
rect 19656 28256 19720 28260
rect 19736 28316 19800 28320
rect 19736 28260 19740 28316
rect 19740 28260 19796 28316
rect 19796 28260 19800 28316
rect 19736 28256 19800 28260
rect 19816 28316 19880 28320
rect 19816 28260 19820 28316
rect 19820 28260 19876 28316
rect 19876 28260 19880 28316
rect 19816 28256 19880 28260
rect 50296 28316 50360 28320
rect 50296 28260 50300 28316
rect 50300 28260 50356 28316
rect 50356 28260 50360 28316
rect 50296 28256 50360 28260
rect 50376 28316 50440 28320
rect 50376 28260 50380 28316
rect 50380 28260 50436 28316
rect 50436 28260 50440 28316
rect 50376 28256 50440 28260
rect 50456 28316 50520 28320
rect 50456 28260 50460 28316
rect 50460 28260 50516 28316
rect 50516 28260 50520 28316
rect 50456 28256 50520 28260
rect 50536 28316 50600 28320
rect 50536 28260 50540 28316
rect 50540 28260 50596 28316
rect 50596 28260 50600 28316
rect 50536 28256 50600 28260
rect 4216 27772 4280 27776
rect 4216 27716 4220 27772
rect 4220 27716 4276 27772
rect 4276 27716 4280 27772
rect 4216 27712 4280 27716
rect 4296 27772 4360 27776
rect 4296 27716 4300 27772
rect 4300 27716 4356 27772
rect 4356 27716 4360 27772
rect 4296 27712 4360 27716
rect 4376 27772 4440 27776
rect 4376 27716 4380 27772
rect 4380 27716 4436 27772
rect 4436 27716 4440 27772
rect 4376 27712 4440 27716
rect 4456 27772 4520 27776
rect 4456 27716 4460 27772
rect 4460 27716 4516 27772
rect 4516 27716 4520 27772
rect 4456 27712 4520 27716
rect 34936 27772 35000 27776
rect 34936 27716 34940 27772
rect 34940 27716 34996 27772
rect 34996 27716 35000 27772
rect 34936 27712 35000 27716
rect 35016 27772 35080 27776
rect 35016 27716 35020 27772
rect 35020 27716 35076 27772
rect 35076 27716 35080 27772
rect 35016 27712 35080 27716
rect 35096 27772 35160 27776
rect 35096 27716 35100 27772
rect 35100 27716 35156 27772
rect 35156 27716 35160 27772
rect 35096 27712 35160 27716
rect 35176 27772 35240 27776
rect 35176 27716 35180 27772
rect 35180 27716 35236 27772
rect 35236 27716 35240 27772
rect 35176 27712 35240 27716
rect 19576 27228 19640 27232
rect 19576 27172 19580 27228
rect 19580 27172 19636 27228
rect 19636 27172 19640 27228
rect 19576 27168 19640 27172
rect 19656 27228 19720 27232
rect 19656 27172 19660 27228
rect 19660 27172 19716 27228
rect 19716 27172 19720 27228
rect 19656 27168 19720 27172
rect 19736 27228 19800 27232
rect 19736 27172 19740 27228
rect 19740 27172 19796 27228
rect 19796 27172 19800 27228
rect 19736 27168 19800 27172
rect 19816 27228 19880 27232
rect 19816 27172 19820 27228
rect 19820 27172 19876 27228
rect 19876 27172 19880 27228
rect 19816 27168 19880 27172
rect 50296 27228 50360 27232
rect 50296 27172 50300 27228
rect 50300 27172 50356 27228
rect 50356 27172 50360 27228
rect 50296 27168 50360 27172
rect 50376 27228 50440 27232
rect 50376 27172 50380 27228
rect 50380 27172 50436 27228
rect 50436 27172 50440 27228
rect 50376 27168 50440 27172
rect 50456 27228 50520 27232
rect 50456 27172 50460 27228
rect 50460 27172 50516 27228
rect 50516 27172 50520 27228
rect 50456 27168 50520 27172
rect 50536 27228 50600 27232
rect 50536 27172 50540 27228
rect 50540 27172 50596 27228
rect 50596 27172 50600 27228
rect 50536 27168 50600 27172
rect 4216 26684 4280 26688
rect 4216 26628 4220 26684
rect 4220 26628 4276 26684
rect 4276 26628 4280 26684
rect 4216 26624 4280 26628
rect 4296 26684 4360 26688
rect 4296 26628 4300 26684
rect 4300 26628 4356 26684
rect 4356 26628 4360 26684
rect 4296 26624 4360 26628
rect 4376 26684 4440 26688
rect 4376 26628 4380 26684
rect 4380 26628 4436 26684
rect 4436 26628 4440 26684
rect 4376 26624 4440 26628
rect 4456 26684 4520 26688
rect 4456 26628 4460 26684
rect 4460 26628 4516 26684
rect 4516 26628 4520 26684
rect 4456 26624 4520 26628
rect 34936 26684 35000 26688
rect 34936 26628 34940 26684
rect 34940 26628 34996 26684
rect 34996 26628 35000 26684
rect 34936 26624 35000 26628
rect 35016 26684 35080 26688
rect 35016 26628 35020 26684
rect 35020 26628 35076 26684
rect 35076 26628 35080 26684
rect 35016 26624 35080 26628
rect 35096 26684 35160 26688
rect 35096 26628 35100 26684
rect 35100 26628 35156 26684
rect 35156 26628 35160 26684
rect 35096 26624 35160 26628
rect 35176 26684 35240 26688
rect 35176 26628 35180 26684
rect 35180 26628 35236 26684
rect 35236 26628 35240 26684
rect 35176 26624 35240 26628
rect 19576 26140 19640 26144
rect 19576 26084 19580 26140
rect 19580 26084 19636 26140
rect 19636 26084 19640 26140
rect 19576 26080 19640 26084
rect 19656 26140 19720 26144
rect 19656 26084 19660 26140
rect 19660 26084 19716 26140
rect 19716 26084 19720 26140
rect 19656 26080 19720 26084
rect 19736 26140 19800 26144
rect 19736 26084 19740 26140
rect 19740 26084 19796 26140
rect 19796 26084 19800 26140
rect 19736 26080 19800 26084
rect 19816 26140 19880 26144
rect 19816 26084 19820 26140
rect 19820 26084 19876 26140
rect 19876 26084 19880 26140
rect 19816 26080 19880 26084
rect 50296 26140 50360 26144
rect 50296 26084 50300 26140
rect 50300 26084 50356 26140
rect 50356 26084 50360 26140
rect 50296 26080 50360 26084
rect 50376 26140 50440 26144
rect 50376 26084 50380 26140
rect 50380 26084 50436 26140
rect 50436 26084 50440 26140
rect 50376 26080 50440 26084
rect 50456 26140 50520 26144
rect 50456 26084 50460 26140
rect 50460 26084 50516 26140
rect 50516 26084 50520 26140
rect 50456 26080 50520 26084
rect 50536 26140 50600 26144
rect 50536 26084 50540 26140
rect 50540 26084 50596 26140
rect 50596 26084 50600 26140
rect 50536 26080 50600 26084
rect 4216 25596 4280 25600
rect 4216 25540 4220 25596
rect 4220 25540 4276 25596
rect 4276 25540 4280 25596
rect 4216 25536 4280 25540
rect 4296 25596 4360 25600
rect 4296 25540 4300 25596
rect 4300 25540 4356 25596
rect 4356 25540 4360 25596
rect 4296 25536 4360 25540
rect 4376 25596 4440 25600
rect 4376 25540 4380 25596
rect 4380 25540 4436 25596
rect 4436 25540 4440 25596
rect 4376 25536 4440 25540
rect 4456 25596 4520 25600
rect 4456 25540 4460 25596
rect 4460 25540 4516 25596
rect 4516 25540 4520 25596
rect 4456 25536 4520 25540
rect 34936 25596 35000 25600
rect 34936 25540 34940 25596
rect 34940 25540 34996 25596
rect 34996 25540 35000 25596
rect 34936 25536 35000 25540
rect 35016 25596 35080 25600
rect 35016 25540 35020 25596
rect 35020 25540 35076 25596
rect 35076 25540 35080 25596
rect 35016 25536 35080 25540
rect 35096 25596 35160 25600
rect 35096 25540 35100 25596
rect 35100 25540 35156 25596
rect 35156 25540 35160 25596
rect 35096 25536 35160 25540
rect 35176 25596 35240 25600
rect 35176 25540 35180 25596
rect 35180 25540 35236 25596
rect 35236 25540 35240 25596
rect 35176 25536 35240 25540
rect 19576 25052 19640 25056
rect 19576 24996 19580 25052
rect 19580 24996 19636 25052
rect 19636 24996 19640 25052
rect 19576 24992 19640 24996
rect 19656 25052 19720 25056
rect 19656 24996 19660 25052
rect 19660 24996 19716 25052
rect 19716 24996 19720 25052
rect 19656 24992 19720 24996
rect 19736 25052 19800 25056
rect 19736 24996 19740 25052
rect 19740 24996 19796 25052
rect 19796 24996 19800 25052
rect 19736 24992 19800 24996
rect 19816 25052 19880 25056
rect 19816 24996 19820 25052
rect 19820 24996 19876 25052
rect 19876 24996 19880 25052
rect 19816 24992 19880 24996
rect 50296 25052 50360 25056
rect 50296 24996 50300 25052
rect 50300 24996 50356 25052
rect 50356 24996 50360 25052
rect 50296 24992 50360 24996
rect 50376 25052 50440 25056
rect 50376 24996 50380 25052
rect 50380 24996 50436 25052
rect 50436 24996 50440 25052
rect 50376 24992 50440 24996
rect 50456 25052 50520 25056
rect 50456 24996 50460 25052
rect 50460 24996 50516 25052
rect 50516 24996 50520 25052
rect 50456 24992 50520 24996
rect 50536 25052 50600 25056
rect 50536 24996 50540 25052
rect 50540 24996 50596 25052
rect 50596 24996 50600 25052
rect 50536 24992 50600 24996
rect 4216 24508 4280 24512
rect 4216 24452 4220 24508
rect 4220 24452 4276 24508
rect 4276 24452 4280 24508
rect 4216 24448 4280 24452
rect 4296 24508 4360 24512
rect 4296 24452 4300 24508
rect 4300 24452 4356 24508
rect 4356 24452 4360 24508
rect 4296 24448 4360 24452
rect 4376 24508 4440 24512
rect 4376 24452 4380 24508
rect 4380 24452 4436 24508
rect 4436 24452 4440 24508
rect 4376 24448 4440 24452
rect 4456 24508 4520 24512
rect 4456 24452 4460 24508
rect 4460 24452 4516 24508
rect 4516 24452 4520 24508
rect 4456 24448 4520 24452
rect 34936 24508 35000 24512
rect 34936 24452 34940 24508
rect 34940 24452 34996 24508
rect 34996 24452 35000 24508
rect 34936 24448 35000 24452
rect 35016 24508 35080 24512
rect 35016 24452 35020 24508
rect 35020 24452 35076 24508
rect 35076 24452 35080 24508
rect 35016 24448 35080 24452
rect 35096 24508 35160 24512
rect 35096 24452 35100 24508
rect 35100 24452 35156 24508
rect 35156 24452 35160 24508
rect 35096 24448 35160 24452
rect 35176 24508 35240 24512
rect 35176 24452 35180 24508
rect 35180 24452 35236 24508
rect 35236 24452 35240 24508
rect 35176 24448 35240 24452
rect 19576 23964 19640 23968
rect 19576 23908 19580 23964
rect 19580 23908 19636 23964
rect 19636 23908 19640 23964
rect 19576 23904 19640 23908
rect 19656 23964 19720 23968
rect 19656 23908 19660 23964
rect 19660 23908 19716 23964
rect 19716 23908 19720 23964
rect 19656 23904 19720 23908
rect 19736 23964 19800 23968
rect 19736 23908 19740 23964
rect 19740 23908 19796 23964
rect 19796 23908 19800 23964
rect 19736 23904 19800 23908
rect 19816 23964 19880 23968
rect 19816 23908 19820 23964
rect 19820 23908 19876 23964
rect 19876 23908 19880 23964
rect 19816 23904 19880 23908
rect 50296 23964 50360 23968
rect 50296 23908 50300 23964
rect 50300 23908 50356 23964
rect 50356 23908 50360 23964
rect 50296 23904 50360 23908
rect 50376 23964 50440 23968
rect 50376 23908 50380 23964
rect 50380 23908 50436 23964
rect 50436 23908 50440 23964
rect 50376 23904 50440 23908
rect 50456 23964 50520 23968
rect 50456 23908 50460 23964
rect 50460 23908 50516 23964
rect 50516 23908 50520 23964
rect 50456 23904 50520 23908
rect 50536 23964 50600 23968
rect 50536 23908 50540 23964
rect 50540 23908 50596 23964
rect 50596 23908 50600 23964
rect 50536 23904 50600 23908
rect 4216 23420 4280 23424
rect 4216 23364 4220 23420
rect 4220 23364 4276 23420
rect 4276 23364 4280 23420
rect 4216 23360 4280 23364
rect 4296 23420 4360 23424
rect 4296 23364 4300 23420
rect 4300 23364 4356 23420
rect 4356 23364 4360 23420
rect 4296 23360 4360 23364
rect 4376 23420 4440 23424
rect 4376 23364 4380 23420
rect 4380 23364 4436 23420
rect 4436 23364 4440 23420
rect 4376 23360 4440 23364
rect 4456 23420 4520 23424
rect 4456 23364 4460 23420
rect 4460 23364 4516 23420
rect 4516 23364 4520 23420
rect 4456 23360 4520 23364
rect 34936 23420 35000 23424
rect 34936 23364 34940 23420
rect 34940 23364 34996 23420
rect 34996 23364 35000 23420
rect 34936 23360 35000 23364
rect 35016 23420 35080 23424
rect 35016 23364 35020 23420
rect 35020 23364 35076 23420
rect 35076 23364 35080 23420
rect 35016 23360 35080 23364
rect 35096 23420 35160 23424
rect 35096 23364 35100 23420
rect 35100 23364 35156 23420
rect 35156 23364 35160 23420
rect 35096 23360 35160 23364
rect 35176 23420 35240 23424
rect 35176 23364 35180 23420
rect 35180 23364 35236 23420
rect 35236 23364 35240 23420
rect 35176 23360 35240 23364
rect 19576 22876 19640 22880
rect 19576 22820 19580 22876
rect 19580 22820 19636 22876
rect 19636 22820 19640 22876
rect 19576 22816 19640 22820
rect 19656 22876 19720 22880
rect 19656 22820 19660 22876
rect 19660 22820 19716 22876
rect 19716 22820 19720 22876
rect 19656 22816 19720 22820
rect 19736 22876 19800 22880
rect 19736 22820 19740 22876
rect 19740 22820 19796 22876
rect 19796 22820 19800 22876
rect 19736 22816 19800 22820
rect 19816 22876 19880 22880
rect 19816 22820 19820 22876
rect 19820 22820 19876 22876
rect 19876 22820 19880 22876
rect 19816 22816 19880 22820
rect 50296 22876 50360 22880
rect 50296 22820 50300 22876
rect 50300 22820 50356 22876
rect 50356 22820 50360 22876
rect 50296 22816 50360 22820
rect 50376 22876 50440 22880
rect 50376 22820 50380 22876
rect 50380 22820 50436 22876
rect 50436 22820 50440 22876
rect 50376 22816 50440 22820
rect 50456 22876 50520 22880
rect 50456 22820 50460 22876
rect 50460 22820 50516 22876
rect 50516 22820 50520 22876
rect 50456 22816 50520 22820
rect 50536 22876 50600 22880
rect 50536 22820 50540 22876
rect 50540 22820 50596 22876
rect 50596 22820 50600 22876
rect 50536 22816 50600 22820
rect 4216 22332 4280 22336
rect 4216 22276 4220 22332
rect 4220 22276 4276 22332
rect 4276 22276 4280 22332
rect 4216 22272 4280 22276
rect 4296 22332 4360 22336
rect 4296 22276 4300 22332
rect 4300 22276 4356 22332
rect 4356 22276 4360 22332
rect 4296 22272 4360 22276
rect 4376 22332 4440 22336
rect 4376 22276 4380 22332
rect 4380 22276 4436 22332
rect 4436 22276 4440 22332
rect 4376 22272 4440 22276
rect 4456 22332 4520 22336
rect 4456 22276 4460 22332
rect 4460 22276 4516 22332
rect 4516 22276 4520 22332
rect 4456 22272 4520 22276
rect 34936 22332 35000 22336
rect 34936 22276 34940 22332
rect 34940 22276 34996 22332
rect 34996 22276 35000 22332
rect 34936 22272 35000 22276
rect 35016 22332 35080 22336
rect 35016 22276 35020 22332
rect 35020 22276 35076 22332
rect 35076 22276 35080 22332
rect 35016 22272 35080 22276
rect 35096 22332 35160 22336
rect 35096 22276 35100 22332
rect 35100 22276 35156 22332
rect 35156 22276 35160 22332
rect 35096 22272 35160 22276
rect 35176 22332 35240 22336
rect 35176 22276 35180 22332
rect 35180 22276 35236 22332
rect 35236 22276 35240 22332
rect 35176 22272 35240 22276
rect 19576 21788 19640 21792
rect 19576 21732 19580 21788
rect 19580 21732 19636 21788
rect 19636 21732 19640 21788
rect 19576 21728 19640 21732
rect 19656 21788 19720 21792
rect 19656 21732 19660 21788
rect 19660 21732 19716 21788
rect 19716 21732 19720 21788
rect 19656 21728 19720 21732
rect 19736 21788 19800 21792
rect 19736 21732 19740 21788
rect 19740 21732 19796 21788
rect 19796 21732 19800 21788
rect 19736 21728 19800 21732
rect 19816 21788 19880 21792
rect 19816 21732 19820 21788
rect 19820 21732 19876 21788
rect 19876 21732 19880 21788
rect 19816 21728 19880 21732
rect 50296 21788 50360 21792
rect 50296 21732 50300 21788
rect 50300 21732 50356 21788
rect 50356 21732 50360 21788
rect 50296 21728 50360 21732
rect 50376 21788 50440 21792
rect 50376 21732 50380 21788
rect 50380 21732 50436 21788
rect 50436 21732 50440 21788
rect 50376 21728 50440 21732
rect 50456 21788 50520 21792
rect 50456 21732 50460 21788
rect 50460 21732 50516 21788
rect 50516 21732 50520 21788
rect 50456 21728 50520 21732
rect 50536 21788 50600 21792
rect 50536 21732 50540 21788
rect 50540 21732 50596 21788
rect 50596 21732 50600 21788
rect 50536 21728 50600 21732
rect 4216 21244 4280 21248
rect 4216 21188 4220 21244
rect 4220 21188 4276 21244
rect 4276 21188 4280 21244
rect 4216 21184 4280 21188
rect 4296 21244 4360 21248
rect 4296 21188 4300 21244
rect 4300 21188 4356 21244
rect 4356 21188 4360 21244
rect 4296 21184 4360 21188
rect 4376 21244 4440 21248
rect 4376 21188 4380 21244
rect 4380 21188 4436 21244
rect 4436 21188 4440 21244
rect 4376 21184 4440 21188
rect 4456 21244 4520 21248
rect 4456 21188 4460 21244
rect 4460 21188 4516 21244
rect 4516 21188 4520 21244
rect 4456 21184 4520 21188
rect 34936 21244 35000 21248
rect 34936 21188 34940 21244
rect 34940 21188 34996 21244
rect 34996 21188 35000 21244
rect 34936 21184 35000 21188
rect 35016 21244 35080 21248
rect 35016 21188 35020 21244
rect 35020 21188 35076 21244
rect 35076 21188 35080 21244
rect 35016 21184 35080 21188
rect 35096 21244 35160 21248
rect 35096 21188 35100 21244
rect 35100 21188 35156 21244
rect 35156 21188 35160 21244
rect 35096 21184 35160 21188
rect 35176 21244 35240 21248
rect 35176 21188 35180 21244
rect 35180 21188 35236 21244
rect 35236 21188 35240 21244
rect 35176 21184 35240 21188
rect 19576 20700 19640 20704
rect 19576 20644 19580 20700
rect 19580 20644 19636 20700
rect 19636 20644 19640 20700
rect 19576 20640 19640 20644
rect 19656 20700 19720 20704
rect 19656 20644 19660 20700
rect 19660 20644 19716 20700
rect 19716 20644 19720 20700
rect 19656 20640 19720 20644
rect 19736 20700 19800 20704
rect 19736 20644 19740 20700
rect 19740 20644 19796 20700
rect 19796 20644 19800 20700
rect 19736 20640 19800 20644
rect 19816 20700 19880 20704
rect 19816 20644 19820 20700
rect 19820 20644 19876 20700
rect 19876 20644 19880 20700
rect 19816 20640 19880 20644
rect 50296 20700 50360 20704
rect 50296 20644 50300 20700
rect 50300 20644 50356 20700
rect 50356 20644 50360 20700
rect 50296 20640 50360 20644
rect 50376 20700 50440 20704
rect 50376 20644 50380 20700
rect 50380 20644 50436 20700
rect 50436 20644 50440 20700
rect 50376 20640 50440 20644
rect 50456 20700 50520 20704
rect 50456 20644 50460 20700
rect 50460 20644 50516 20700
rect 50516 20644 50520 20700
rect 50456 20640 50520 20644
rect 50536 20700 50600 20704
rect 50536 20644 50540 20700
rect 50540 20644 50596 20700
rect 50596 20644 50600 20700
rect 50536 20640 50600 20644
rect 4216 20156 4280 20160
rect 4216 20100 4220 20156
rect 4220 20100 4276 20156
rect 4276 20100 4280 20156
rect 4216 20096 4280 20100
rect 4296 20156 4360 20160
rect 4296 20100 4300 20156
rect 4300 20100 4356 20156
rect 4356 20100 4360 20156
rect 4296 20096 4360 20100
rect 4376 20156 4440 20160
rect 4376 20100 4380 20156
rect 4380 20100 4436 20156
rect 4436 20100 4440 20156
rect 4376 20096 4440 20100
rect 4456 20156 4520 20160
rect 4456 20100 4460 20156
rect 4460 20100 4516 20156
rect 4516 20100 4520 20156
rect 4456 20096 4520 20100
rect 34936 20156 35000 20160
rect 34936 20100 34940 20156
rect 34940 20100 34996 20156
rect 34996 20100 35000 20156
rect 34936 20096 35000 20100
rect 35016 20156 35080 20160
rect 35016 20100 35020 20156
rect 35020 20100 35076 20156
rect 35076 20100 35080 20156
rect 35016 20096 35080 20100
rect 35096 20156 35160 20160
rect 35096 20100 35100 20156
rect 35100 20100 35156 20156
rect 35156 20100 35160 20156
rect 35096 20096 35160 20100
rect 35176 20156 35240 20160
rect 35176 20100 35180 20156
rect 35180 20100 35236 20156
rect 35236 20100 35240 20156
rect 35176 20096 35240 20100
rect 19576 19612 19640 19616
rect 19576 19556 19580 19612
rect 19580 19556 19636 19612
rect 19636 19556 19640 19612
rect 19576 19552 19640 19556
rect 19656 19612 19720 19616
rect 19656 19556 19660 19612
rect 19660 19556 19716 19612
rect 19716 19556 19720 19612
rect 19656 19552 19720 19556
rect 19736 19612 19800 19616
rect 19736 19556 19740 19612
rect 19740 19556 19796 19612
rect 19796 19556 19800 19612
rect 19736 19552 19800 19556
rect 19816 19612 19880 19616
rect 19816 19556 19820 19612
rect 19820 19556 19876 19612
rect 19876 19556 19880 19612
rect 19816 19552 19880 19556
rect 50296 19612 50360 19616
rect 50296 19556 50300 19612
rect 50300 19556 50356 19612
rect 50356 19556 50360 19612
rect 50296 19552 50360 19556
rect 50376 19612 50440 19616
rect 50376 19556 50380 19612
rect 50380 19556 50436 19612
rect 50436 19556 50440 19612
rect 50376 19552 50440 19556
rect 50456 19612 50520 19616
rect 50456 19556 50460 19612
rect 50460 19556 50516 19612
rect 50516 19556 50520 19612
rect 50456 19552 50520 19556
rect 50536 19612 50600 19616
rect 50536 19556 50540 19612
rect 50540 19556 50596 19612
rect 50596 19556 50600 19612
rect 50536 19552 50600 19556
rect 4216 19068 4280 19072
rect 4216 19012 4220 19068
rect 4220 19012 4276 19068
rect 4276 19012 4280 19068
rect 4216 19008 4280 19012
rect 4296 19068 4360 19072
rect 4296 19012 4300 19068
rect 4300 19012 4356 19068
rect 4356 19012 4360 19068
rect 4296 19008 4360 19012
rect 4376 19068 4440 19072
rect 4376 19012 4380 19068
rect 4380 19012 4436 19068
rect 4436 19012 4440 19068
rect 4376 19008 4440 19012
rect 4456 19068 4520 19072
rect 4456 19012 4460 19068
rect 4460 19012 4516 19068
rect 4516 19012 4520 19068
rect 4456 19008 4520 19012
rect 34936 19068 35000 19072
rect 34936 19012 34940 19068
rect 34940 19012 34996 19068
rect 34996 19012 35000 19068
rect 34936 19008 35000 19012
rect 35016 19068 35080 19072
rect 35016 19012 35020 19068
rect 35020 19012 35076 19068
rect 35076 19012 35080 19068
rect 35016 19008 35080 19012
rect 35096 19068 35160 19072
rect 35096 19012 35100 19068
rect 35100 19012 35156 19068
rect 35156 19012 35160 19068
rect 35096 19008 35160 19012
rect 35176 19068 35240 19072
rect 35176 19012 35180 19068
rect 35180 19012 35236 19068
rect 35236 19012 35240 19068
rect 35176 19008 35240 19012
rect 19576 18524 19640 18528
rect 19576 18468 19580 18524
rect 19580 18468 19636 18524
rect 19636 18468 19640 18524
rect 19576 18464 19640 18468
rect 19656 18524 19720 18528
rect 19656 18468 19660 18524
rect 19660 18468 19716 18524
rect 19716 18468 19720 18524
rect 19656 18464 19720 18468
rect 19736 18524 19800 18528
rect 19736 18468 19740 18524
rect 19740 18468 19796 18524
rect 19796 18468 19800 18524
rect 19736 18464 19800 18468
rect 19816 18524 19880 18528
rect 19816 18468 19820 18524
rect 19820 18468 19876 18524
rect 19876 18468 19880 18524
rect 19816 18464 19880 18468
rect 50296 18524 50360 18528
rect 50296 18468 50300 18524
rect 50300 18468 50356 18524
rect 50356 18468 50360 18524
rect 50296 18464 50360 18468
rect 50376 18524 50440 18528
rect 50376 18468 50380 18524
rect 50380 18468 50436 18524
rect 50436 18468 50440 18524
rect 50376 18464 50440 18468
rect 50456 18524 50520 18528
rect 50456 18468 50460 18524
rect 50460 18468 50516 18524
rect 50516 18468 50520 18524
rect 50456 18464 50520 18468
rect 50536 18524 50600 18528
rect 50536 18468 50540 18524
rect 50540 18468 50596 18524
rect 50596 18468 50600 18524
rect 50536 18464 50600 18468
rect 4216 17980 4280 17984
rect 4216 17924 4220 17980
rect 4220 17924 4276 17980
rect 4276 17924 4280 17980
rect 4216 17920 4280 17924
rect 4296 17980 4360 17984
rect 4296 17924 4300 17980
rect 4300 17924 4356 17980
rect 4356 17924 4360 17980
rect 4296 17920 4360 17924
rect 4376 17980 4440 17984
rect 4376 17924 4380 17980
rect 4380 17924 4436 17980
rect 4436 17924 4440 17980
rect 4376 17920 4440 17924
rect 4456 17980 4520 17984
rect 4456 17924 4460 17980
rect 4460 17924 4516 17980
rect 4516 17924 4520 17980
rect 4456 17920 4520 17924
rect 34936 17980 35000 17984
rect 34936 17924 34940 17980
rect 34940 17924 34996 17980
rect 34996 17924 35000 17980
rect 34936 17920 35000 17924
rect 35016 17980 35080 17984
rect 35016 17924 35020 17980
rect 35020 17924 35076 17980
rect 35076 17924 35080 17980
rect 35016 17920 35080 17924
rect 35096 17980 35160 17984
rect 35096 17924 35100 17980
rect 35100 17924 35156 17980
rect 35156 17924 35160 17980
rect 35096 17920 35160 17924
rect 35176 17980 35240 17984
rect 35176 17924 35180 17980
rect 35180 17924 35236 17980
rect 35236 17924 35240 17980
rect 35176 17920 35240 17924
rect 19576 17436 19640 17440
rect 19576 17380 19580 17436
rect 19580 17380 19636 17436
rect 19636 17380 19640 17436
rect 19576 17376 19640 17380
rect 19656 17436 19720 17440
rect 19656 17380 19660 17436
rect 19660 17380 19716 17436
rect 19716 17380 19720 17436
rect 19656 17376 19720 17380
rect 19736 17436 19800 17440
rect 19736 17380 19740 17436
rect 19740 17380 19796 17436
rect 19796 17380 19800 17436
rect 19736 17376 19800 17380
rect 19816 17436 19880 17440
rect 19816 17380 19820 17436
rect 19820 17380 19876 17436
rect 19876 17380 19880 17436
rect 19816 17376 19880 17380
rect 50296 17436 50360 17440
rect 50296 17380 50300 17436
rect 50300 17380 50356 17436
rect 50356 17380 50360 17436
rect 50296 17376 50360 17380
rect 50376 17436 50440 17440
rect 50376 17380 50380 17436
rect 50380 17380 50436 17436
rect 50436 17380 50440 17436
rect 50376 17376 50440 17380
rect 50456 17436 50520 17440
rect 50456 17380 50460 17436
rect 50460 17380 50516 17436
rect 50516 17380 50520 17436
rect 50456 17376 50520 17380
rect 50536 17436 50600 17440
rect 50536 17380 50540 17436
rect 50540 17380 50596 17436
rect 50596 17380 50600 17436
rect 50536 17376 50600 17380
rect 4216 16892 4280 16896
rect 4216 16836 4220 16892
rect 4220 16836 4276 16892
rect 4276 16836 4280 16892
rect 4216 16832 4280 16836
rect 4296 16892 4360 16896
rect 4296 16836 4300 16892
rect 4300 16836 4356 16892
rect 4356 16836 4360 16892
rect 4296 16832 4360 16836
rect 4376 16892 4440 16896
rect 4376 16836 4380 16892
rect 4380 16836 4436 16892
rect 4436 16836 4440 16892
rect 4376 16832 4440 16836
rect 4456 16892 4520 16896
rect 4456 16836 4460 16892
rect 4460 16836 4516 16892
rect 4516 16836 4520 16892
rect 4456 16832 4520 16836
rect 34936 16892 35000 16896
rect 34936 16836 34940 16892
rect 34940 16836 34996 16892
rect 34996 16836 35000 16892
rect 34936 16832 35000 16836
rect 35016 16892 35080 16896
rect 35016 16836 35020 16892
rect 35020 16836 35076 16892
rect 35076 16836 35080 16892
rect 35016 16832 35080 16836
rect 35096 16892 35160 16896
rect 35096 16836 35100 16892
rect 35100 16836 35156 16892
rect 35156 16836 35160 16892
rect 35096 16832 35160 16836
rect 35176 16892 35240 16896
rect 35176 16836 35180 16892
rect 35180 16836 35236 16892
rect 35236 16836 35240 16892
rect 35176 16832 35240 16836
rect 19576 16348 19640 16352
rect 19576 16292 19580 16348
rect 19580 16292 19636 16348
rect 19636 16292 19640 16348
rect 19576 16288 19640 16292
rect 19656 16348 19720 16352
rect 19656 16292 19660 16348
rect 19660 16292 19716 16348
rect 19716 16292 19720 16348
rect 19656 16288 19720 16292
rect 19736 16348 19800 16352
rect 19736 16292 19740 16348
rect 19740 16292 19796 16348
rect 19796 16292 19800 16348
rect 19736 16288 19800 16292
rect 19816 16348 19880 16352
rect 19816 16292 19820 16348
rect 19820 16292 19876 16348
rect 19876 16292 19880 16348
rect 19816 16288 19880 16292
rect 50296 16348 50360 16352
rect 50296 16292 50300 16348
rect 50300 16292 50356 16348
rect 50356 16292 50360 16348
rect 50296 16288 50360 16292
rect 50376 16348 50440 16352
rect 50376 16292 50380 16348
rect 50380 16292 50436 16348
rect 50436 16292 50440 16348
rect 50376 16288 50440 16292
rect 50456 16348 50520 16352
rect 50456 16292 50460 16348
rect 50460 16292 50516 16348
rect 50516 16292 50520 16348
rect 50456 16288 50520 16292
rect 50536 16348 50600 16352
rect 50536 16292 50540 16348
rect 50540 16292 50596 16348
rect 50596 16292 50600 16348
rect 50536 16288 50600 16292
rect 4216 15804 4280 15808
rect 4216 15748 4220 15804
rect 4220 15748 4276 15804
rect 4276 15748 4280 15804
rect 4216 15744 4280 15748
rect 4296 15804 4360 15808
rect 4296 15748 4300 15804
rect 4300 15748 4356 15804
rect 4356 15748 4360 15804
rect 4296 15744 4360 15748
rect 4376 15804 4440 15808
rect 4376 15748 4380 15804
rect 4380 15748 4436 15804
rect 4436 15748 4440 15804
rect 4376 15744 4440 15748
rect 4456 15804 4520 15808
rect 4456 15748 4460 15804
rect 4460 15748 4516 15804
rect 4516 15748 4520 15804
rect 4456 15744 4520 15748
rect 34936 15804 35000 15808
rect 34936 15748 34940 15804
rect 34940 15748 34996 15804
rect 34996 15748 35000 15804
rect 34936 15744 35000 15748
rect 35016 15804 35080 15808
rect 35016 15748 35020 15804
rect 35020 15748 35076 15804
rect 35076 15748 35080 15804
rect 35016 15744 35080 15748
rect 35096 15804 35160 15808
rect 35096 15748 35100 15804
rect 35100 15748 35156 15804
rect 35156 15748 35160 15804
rect 35096 15744 35160 15748
rect 35176 15804 35240 15808
rect 35176 15748 35180 15804
rect 35180 15748 35236 15804
rect 35236 15748 35240 15804
rect 35176 15744 35240 15748
rect 19576 15260 19640 15264
rect 19576 15204 19580 15260
rect 19580 15204 19636 15260
rect 19636 15204 19640 15260
rect 19576 15200 19640 15204
rect 19656 15260 19720 15264
rect 19656 15204 19660 15260
rect 19660 15204 19716 15260
rect 19716 15204 19720 15260
rect 19656 15200 19720 15204
rect 19736 15260 19800 15264
rect 19736 15204 19740 15260
rect 19740 15204 19796 15260
rect 19796 15204 19800 15260
rect 19736 15200 19800 15204
rect 19816 15260 19880 15264
rect 19816 15204 19820 15260
rect 19820 15204 19876 15260
rect 19876 15204 19880 15260
rect 19816 15200 19880 15204
rect 50296 15260 50360 15264
rect 50296 15204 50300 15260
rect 50300 15204 50356 15260
rect 50356 15204 50360 15260
rect 50296 15200 50360 15204
rect 50376 15260 50440 15264
rect 50376 15204 50380 15260
rect 50380 15204 50436 15260
rect 50436 15204 50440 15260
rect 50376 15200 50440 15204
rect 50456 15260 50520 15264
rect 50456 15204 50460 15260
rect 50460 15204 50516 15260
rect 50516 15204 50520 15260
rect 50456 15200 50520 15204
rect 50536 15260 50600 15264
rect 50536 15204 50540 15260
rect 50540 15204 50596 15260
rect 50596 15204 50600 15260
rect 50536 15200 50600 15204
rect 4216 14716 4280 14720
rect 4216 14660 4220 14716
rect 4220 14660 4276 14716
rect 4276 14660 4280 14716
rect 4216 14656 4280 14660
rect 4296 14716 4360 14720
rect 4296 14660 4300 14716
rect 4300 14660 4356 14716
rect 4356 14660 4360 14716
rect 4296 14656 4360 14660
rect 4376 14716 4440 14720
rect 4376 14660 4380 14716
rect 4380 14660 4436 14716
rect 4436 14660 4440 14716
rect 4376 14656 4440 14660
rect 4456 14716 4520 14720
rect 4456 14660 4460 14716
rect 4460 14660 4516 14716
rect 4516 14660 4520 14716
rect 4456 14656 4520 14660
rect 34936 14716 35000 14720
rect 34936 14660 34940 14716
rect 34940 14660 34996 14716
rect 34996 14660 35000 14716
rect 34936 14656 35000 14660
rect 35016 14716 35080 14720
rect 35016 14660 35020 14716
rect 35020 14660 35076 14716
rect 35076 14660 35080 14716
rect 35016 14656 35080 14660
rect 35096 14716 35160 14720
rect 35096 14660 35100 14716
rect 35100 14660 35156 14716
rect 35156 14660 35160 14716
rect 35096 14656 35160 14660
rect 35176 14716 35240 14720
rect 35176 14660 35180 14716
rect 35180 14660 35236 14716
rect 35236 14660 35240 14716
rect 35176 14656 35240 14660
rect 19576 14172 19640 14176
rect 19576 14116 19580 14172
rect 19580 14116 19636 14172
rect 19636 14116 19640 14172
rect 19576 14112 19640 14116
rect 19656 14172 19720 14176
rect 19656 14116 19660 14172
rect 19660 14116 19716 14172
rect 19716 14116 19720 14172
rect 19656 14112 19720 14116
rect 19736 14172 19800 14176
rect 19736 14116 19740 14172
rect 19740 14116 19796 14172
rect 19796 14116 19800 14172
rect 19736 14112 19800 14116
rect 19816 14172 19880 14176
rect 19816 14116 19820 14172
rect 19820 14116 19876 14172
rect 19876 14116 19880 14172
rect 19816 14112 19880 14116
rect 50296 14172 50360 14176
rect 50296 14116 50300 14172
rect 50300 14116 50356 14172
rect 50356 14116 50360 14172
rect 50296 14112 50360 14116
rect 50376 14172 50440 14176
rect 50376 14116 50380 14172
rect 50380 14116 50436 14172
rect 50436 14116 50440 14172
rect 50376 14112 50440 14116
rect 50456 14172 50520 14176
rect 50456 14116 50460 14172
rect 50460 14116 50516 14172
rect 50516 14116 50520 14172
rect 50456 14112 50520 14116
rect 50536 14172 50600 14176
rect 50536 14116 50540 14172
rect 50540 14116 50596 14172
rect 50596 14116 50600 14172
rect 50536 14112 50600 14116
rect 4216 13628 4280 13632
rect 4216 13572 4220 13628
rect 4220 13572 4276 13628
rect 4276 13572 4280 13628
rect 4216 13568 4280 13572
rect 4296 13628 4360 13632
rect 4296 13572 4300 13628
rect 4300 13572 4356 13628
rect 4356 13572 4360 13628
rect 4296 13568 4360 13572
rect 4376 13628 4440 13632
rect 4376 13572 4380 13628
rect 4380 13572 4436 13628
rect 4436 13572 4440 13628
rect 4376 13568 4440 13572
rect 4456 13628 4520 13632
rect 4456 13572 4460 13628
rect 4460 13572 4516 13628
rect 4516 13572 4520 13628
rect 4456 13568 4520 13572
rect 34936 13628 35000 13632
rect 34936 13572 34940 13628
rect 34940 13572 34996 13628
rect 34996 13572 35000 13628
rect 34936 13568 35000 13572
rect 35016 13628 35080 13632
rect 35016 13572 35020 13628
rect 35020 13572 35076 13628
rect 35076 13572 35080 13628
rect 35016 13568 35080 13572
rect 35096 13628 35160 13632
rect 35096 13572 35100 13628
rect 35100 13572 35156 13628
rect 35156 13572 35160 13628
rect 35096 13568 35160 13572
rect 35176 13628 35240 13632
rect 35176 13572 35180 13628
rect 35180 13572 35236 13628
rect 35236 13572 35240 13628
rect 35176 13568 35240 13572
rect 19576 13084 19640 13088
rect 19576 13028 19580 13084
rect 19580 13028 19636 13084
rect 19636 13028 19640 13084
rect 19576 13024 19640 13028
rect 19656 13084 19720 13088
rect 19656 13028 19660 13084
rect 19660 13028 19716 13084
rect 19716 13028 19720 13084
rect 19656 13024 19720 13028
rect 19736 13084 19800 13088
rect 19736 13028 19740 13084
rect 19740 13028 19796 13084
rect 19796 13028 19800 13084
rect 19736 13024 19800 13028
rect 19816 13084 19880 13088
rect 19816 13028 19820 13084
rect 19820 13028 19876 13084
rect 19876 13028 19880 13084
rect 19816 13024 19880 13028
rect 50296 13084 50360 13088
rect 50296 13028 50300 13084
rect 50300 13028 50356 13084
rect 50356 13028 50360 13084
rect 50296 13024 50360 13028
rect 50376 13084 50440 13088
rect 50376 13028 50380 13084
rect 50380 13028 50436 13084
rect 50436 13028 50440 13084
rect 50376 13024 50440 13028
rect 50456 13084 50520 13088
rect 50456 13028 50460 13084
rect 50460 13028 50516 13084
rect 50516 13028 50520 13084
rect 50456 13024 50520 13028
rect 50536 13084 50600 13088
rect 50536 13028 50540 13084
rect 50540 13028 50596 13084
rect 50596 13028 50600 13084
rect 50536 13024 50600 13028
rect 4216 12540 4280 12544
rect 4216 12484 4220 12540
rect 4220 12484 4276 12540
rect 4276 12484 4280 12540
rect 4216 12480 4280 12484
rect 4296 12540 4360 12544
rect 4296 12484 4300 12540
rect 4300 12484 4356 12540
rect 4356 12484 4360 12540
rect 4296 12480 4360 12484
rect 4376 12540 4440 12544
rect 4376 12484 4380 12540
rect 4380 12484 4436 12540
rect 4436 12484 4440 12540
rect 4376 12480 4440 12484
rect 4456 12540 4520 12544
rect 4456 12484 4460 12540
rect 4460 12484 4516 12540
rect 4516 12484 4520 12540
rect 4456 12480 4520 12484
rect 34936 12540 35000 12544
rect 34936 12484 34940 12540
rect 34940 12484 34996 12540
rect 34996 12484 35000 12540
rect 34936 12480 35000 12484
rect 35016 12540 35080 12544
rect 35016 12484 35020 12540
rect 35020 12484 35076 12540
rect 35076 12484 35080 12540
rect 35016 12480 35080 12484
rect 35096 12540 35160 12544
rect 35096 12484 35100 12540
rect 35100 12484 35156 12540
rect 35156 12484 35160 12540
rect 35096 12480 35160 12484
rect 35176 12540 35240 12544
rect 35176 12484 35180 12540
rect 35180 12484 35236 12540
rect 35236 12484 35240 12540
rect 35176 12480 35240 12484
rect 19576 11996 19640 12000
rect 19576 11940 19580 11996
rect 19580 11940 19636 11996
rect 19636 11940 19640 11996
rect 19576 11936 19640 11940
rect 19656 11996 19720 12000
rect 19656 11940 19660 11996
rect 19660 11940 19716 11996
rect 19716 11940 19720 11996
rect 19656 11936 19720 11940
rect 19736 11996 19800 12000
rect 19736 11940 19740 11996
rect 19740 11940 19796 11996
rect 19796 11940 19800 11996
rect 19736 11936 19800 11940
rect 19816 11996 19880 12000
rect 19816 11940 19820 11996
rect 19820 11940 19876 11996
rect 19876 11940 19880 11996
rect 19816 11936 19880 11940
rect 50296 11996 50360 12000
rect 50296 11940 50300 11996
rect 50300 11940 50356 11996
rect 50356 11940 50360 11996
rect 50296 11936 50360 11940
rect 50376 11996 50440 12000
rect 50376 11940 50380 11996
rect 50380 11940 50436 11996
rect 50436 11940 50440 11996
rect 50376 11936 50440 11940
rect 50456 11996 50520 12000
rect 50456 11940 50460 11996
rect 50460 11940 50516 11996
rect 50516 11940 50520 11996
rect 50456 11936 50520 11940
rect 50536 11996 50600 12000
rect 50536 11940 50540 11996
rect 50540 11940 50596 11996
rect 50596 11940 50600 11996
rect 50536 11936 50600 11940
rect 4216 11452 4280 11456
rect 4216 11396 4220 11452
rect 4220 11396 4276 11452
rect 4276 11396 4280 11452
rect 4216 11392 4280 11396
rect 4296 11452 4360 11456
rect 4296 11396 4300 11452
rect 4300 11396 4356 11452
rect 4356 11396 4360 11452
rect 4296 11392 4360 11396
rect 4376 11452 4440 11456
rect 4376 11396 4380 11452
rect 4380 11396 4436 11452
rect 4436 11396 4440 11452
rect 4376 11392 4440 11396
rect 4456 11452 4520 11456
rect 4456 11396 4460 11452
rect 4460 11396 4516 11452
rect 4516 11396 4520 11452
rect 4456 11392 4520 11396
rect 34936 11452 35000 11456
rect 34936 11396 34940 11452
rect 34940 11396 34996 11452
rect 34996 11396 35000 11452
rect 34936 11392 35000 11396
rect 35016 11452 35080 11456
rect 35016 11396 35020 11452
rect 35020 11396 35076 11452
rect 35076 11396 35080 11452
rect 35016 11392 35080 11396
rect 35096 11452 35160 11456
rect 35096 11396 35100 11452
rect 35100 11396 35156 11452
rect 35156 11396 35160 11452
rect 35096 11392 35160 11396
rect 35176 11452 35240 11456
rect 35176 11396 35180 11452
rect 35180 11396 35236 11452
rect 35236 11396 35240 11452
rect 35176 11392 35240 11396
rect 19576 10908 19640 10912
rect 19576 10852 19580 10908
rect 19580 10852 19636 10908
rect 19636 10852 19640 10908
rect 19576 10848 19640 10852
rect 19656 10908 19720 10912
rect 19656 10852 19660 10908
rect 19660 10852 19716 10908
rect 19716 10852 19720 10908
rect 19656 10848 19720 10852
rect 19736 10908 19800 10912
rect 19736 10852 19740 10908
rect 19740 10852 19796 10908
rect 19796 10852 19800 10908
rect 19736 10848 19800 10852
rect 19816 10908 19880 10912
rect 19816 10852 19820 10908
rect 19820 10852 19876 10908
rect 19876 10852 19880 10908
rect 19816 10848 19880 10852
rect 50296 10908 50360 10912
rect 50296 10852 50300 10908
rect 50300 10852 50356 10908
rect 50356 10852 50360 10908
rect 50296 10848 50360 10852
rect 50376 10908 50440 10912
rect 50376 10852 50380 10908
rect 50380 10852 50436 10908
rect 50436 10852 50440 10908
rect 50376 10848 50440 10852
rect 50456 10908 50520 10912
rect 50456 10852 50460 10908
rect 50460 10852 50516 10908
rect 50516 10852 50520 10908
rect 50456 10848 50520 10852
rect 50536 10908 50600 10912
rect 50536 10852 50540 10908
rect 50540 10852 50596 10908
rect 50596 10852 50600 10908
rect 50536 10848 50600 10852
rect 4216 10364 4280 10368
rect 4216 10308 4220 10364
rect 4220 10308 4276 10364
rect 4276 10308 4280 10364
rect 4216 10304 4280 10308
rect 4296 10364 4360 10368
rect 4296 10308 4300 10364
rect 4300 10308 4356 10364
rect 4356 10308 4360 10364
rect 4296 10304 4360 10308
rect 4376 10364 4440 10368
rect 4376 10308 4380 10364
rect 4380 10308 4436 10364
rect 4436 10308 4440 10364
rect 4376 10304 4440 10308
rect 4456 10364 4520 10368
rect 4456 10308 4460 10364
rect 4460 10308 4516 10364
rect 4516 10308 4520 10364
rect 4456 10304 4520 10308
rect 34936 10364 35000 10368
rect 34936 10308 34940 10364
rect 34940 10308 34996 10364
rect 34996 10308 35000 10364
rect 34936 10304 35000 10308
rect 35016 10364 35080 10368
rect 35016 10308 35020 10364
rect 35020 10308 35076 10364
rect 35076 10308 35080 10364
rect 35016 10304 35080 10308
rect 35096 10364 35160 10368
rect 35096 10308 35100 10364
rect 35100 10308 35156 10364
rect 35156 10308 35160 10364
rect 35096 10304 35160 10308
rect 35176 10364 35240 10368
rect 35176 10308 35180 10364
rect 35180 10308 35236 10364
rect 35236 10308 35240 10364
rect 35176 10304 35240 10308
rect 19576 9820 19640 9824
rect 19576 9764 19580 9820
rect 19580 9764 19636 9820
rect 19636 9764 19640 9820
rect 19576 9760 19640 9764
rect 19656 9820 19720 9824
rect 19656 9764 19660 9820
rect 19660 9764 19716 9820
rect 19716 9764 19720 9820
rect 19656 9760 19720 9764
rect 19736 9820 19800 9824
rect 19736 9764 19740 9820
rect 19740 9764 19796 9820
rect 19796 9764 19800 9820
rect 19736 9760 19800 9764
rect 19816 9820 19880 9824
rect 19816 9764 19820 9820
rect 19820 9764 19876 9820
rect 19876 9764 19880 9820
rect 19816 9760 19880 9764
rect 50296 9820 50360 9824
rect 50296 9764 50300 9820
rect 50300 9764 50356 9820
rect 50356 9764 50360 9820
rect 50296 9760 50360 9764
rect 50376 9820 50440 9824
rect 50376 9764 50380 9820
rect 50380 9764 50436 9820
rect 50436 9764 50440 9820
rect 50376 9760 50440 9764
rect 50456 9820 50520 9824
rect 50456 9764 50460 9820
rect 50460 9764 50516 9820
rect 50516 9764 50520 9820
rect 50456 9760 50520 9764
rect 50536 9820 50600 9824
rect 50536 9764 50540 9820
rect 50540 9764 50596 9820
rect 50596 9764 50600 9820
rect 50536 9760 50600 9764
rect 4216 9276 4280 9280
rect 4216 9220 4220 9276
rect 4220 9220 4276 9276
rect 4276 9220 4280 9276
rect 4216 9216 4280 9220
rect 4296 9276 4360 9280
rect 4296 9220 4300 9276
rect 4300 9220 4356 9276
rect 4356 9220 4360 9276
rect 4296 9216 4360 9220
rect 4376 9276 4440 9280
rect 4376 9220 4380 9276
rect 4380 9220 4436 9276
rect 4436 9220 4440 9276
rect 4376 9216 4440 9220
rect 4456 9276 4520 9280
rect 4456 9220 4460 9276
rect 4460 9220 4516 9276
rect 4516 9220 4520 9276
rect 4456 9216 4520 9220
rect 34936 9276 35000 9280
rect 34936 9220 34940 9276
rect 34940 9220 34996 9276
rect 34996 9220 35000 9276
rect 34936 9216 35000 9220
rect 35016 9276 35080 9280
rect 35016 9220 35020 9276
rect 35020 9220 35076 9276
rect 35076 9220 35080 9276
rect 35016 9216 35080 9220
rect 35096 9276 35160 9280
rect 35096 9220 35100 9276
rect 35100 9220 35156 9276
rect 35156 9220 35160 9276
rect 35096 9216 35160 9220
rect 35176 9276 35240 9280
rect 35176 9220 35180 9276
rect 35180 9220 35236 9276
rect 35236 9220 35240 9276
rect 35176 9216 35240 9220
rect 19576 8732 19640 8736
rect 19576 8676 19580 8732
rect 19580 8676 19636 8732
rect 19636 8676 19640 8732
rect 19576 8672 19640 8676
rect 19656 8732 19720 8736
rect 19656 8676 19660 8732
rect 19660 8676 19716 8732
rect 19716 8676 19720 8732
rect 19656 8672 19720 8676
rect 19736 8732 19800 8736
rect 19736 8676 19740 8732
rect 19740 8676 19796 8732
rect 19796 8676 19800 8732
rect 19736 8672 19800 8676
rect 19816 8732 19880 8736
rect 19816 8676 19820 8732
rect 19820 8676 19876 8732
rect 19876 8676 19880 8732
rect 19816 8672 19880 8676
rect 50296 8732 50360 8736
rect 50296 8676 50300 8732
rect 50300 8676 50356 8732
rect 50356 8676 50360 8732
rect 50296 8672 50360 8676
rect 50376 8732 50440 8736
rect 50376 8676 50380 8732
rect 50380 8676 50436 8732
rect 50436 8676 50440 8732
rect 50376 8672 50440 8676
rect 50456 8732 50520 8736
rect 50456 8676 50460 8732
rect 50460 8676 50516 8732
rect 50516 8676 50520 8732
rect 50456 8672 50520 8676
rect 50536 8732 50600 8736
rect 50536 8676 50540 8732
rect 50540 8676 50596 8732
rect 50596 8676 50600 8732
rect 50536 8672 50600 8676
rect 4216 8188 4280 8192
rect 4216 8132 4220 8188
rect 4220 8132 4276 8188
rect 4276 8132 4280 8188
rect 4216 8128 4280 8132
rect 4296 8188 4360 8192
rect 4296 8132 4300 8188
rect 4300 8132 4356 8188
rect 4356 8132 4360 8188
rect 4296 8128 4360 8132
rect 4376 8188 4440 8192
rect 4376 8132 4380 8188
rect 4380 8132 4436 8188
rect 4436 8132 4440 8188
rect 4376 8128 4440 8132
rect 4456 8188 4520 8192
rect 4456 8132 4460 8188
rect 4460 8132 4516 8188
rect 4516 8132 4520 8188
rect 4456 8128 4520 8132
rect 34936 8188 35000 8192
rect 34936 8132 34940 8188
rect 34940 8132 34996 8188
rect 34996 8132 35000 8188
rect 34936 8128 35000 8132
rect 35016 8188 35080 8192
rect 35016 8132 35020 8188
rect 35020 8132 35076 8188
rect 35076 8132 35080 8188
rect 35016 8128 35080 8132
rect 35096 8188 35160 8192
rect 35096 8132 35100 8188
rect 35100 8132 35156 8188
rect 35156 8132 35160 8188
rect 35096 8128 35160 8132
rect 35176 8188 35240 8192
rect 35176 8132 35180 8188
rect 35180 8132 35236 8188
rect 35236 8132 35240 8188
rect 35176 8128 35240 8132
rect 19576 7644 19640 7648
rect 19576 7588 19580 7644
rect 19580 7588 19636 7644
rect 19636 7588 19640 7644
rect 19576 7584 19640 7588
rect 19656 7644 19720 7648
rect 19656 7588 19660 7644
rect 19660 7588 19716 7644
rect 19716 7588 19720 7644
rect 19656 7584 19720 7588
rect 19736 7644 19800 7648
rect 19736 7588 19740 7644
rect 19740 7588 19796 7644
rect 19796 7588 19800 7644
rect 19736 7584 19800 7588
rect 19816 7644 19880 7648
rect 19816 7588 19820 7644
rect 19820 7588 19876 7644
rect 19876 7588 19880 7644
rect 19816 7584 19880 7588
rect 50296 7644 50360 7648
rect 50296 7588 50300 7644
rect 50300 7588 50356 7644
rect 50356 7588 50360 7644
rect 50296 7584 50360 7588
rect 50376 7644 50440 7648
rect 50376 7588 50380 7644
rect 50380 7588 50436 7644
rect 50436 7588 50440 7644
rect 50376 7584 50440 7588
rect 50456 7644 50520 7648
rect 50456 7588 50460 7644
rect 50460 7588 50516 7644
rect 50516 7588 50520 7644
rect 50456 7584 50520 7588
rect 50536 7644 50600 7648
rect 50536 7588 50540 7644
rect 50540 7588 50596 7644
rect 50596 7588 50600 7644
rect 50536 7584 50600 7588
rect 4216 7100 4280 7104
rect 4216 7044 4220 7100
rect 4220 7044 4276 7100
rect 4276 7044 4280 7100
rect 4216 7040 4280 7044
rect 4296 7100 4360 7104
rect 4296 7044 4300 7100
rect 4300 7044 4356 7100
rect 4356 7044 4360 7100
rect 4296 7040 4360 7044
rect 4376 7100 4440 7104
rect 4376 7044 4380 7100
rect 4380 7044 4436 7100
rect 4436 7044 4440 7100
rect 4376 7040 4440 7044
rect 4456 7100 4520 7104
rect 4456 7044 4460 7100
rect 4460 7044 4516 7100
rect 4516 7044 4520 7100
rect 4456 7040 4520 7044
rect 34936 7100 35000 7104
rect 34936 7044 34940 7100
rect 34940 7044 34996 7100
rect 34996 7044 35000 7100
rect 34936 7040 35000 7044
rect 35016 7100 35080 7104
rect 35016 7044 35020 7100
rect 35020 7044 35076 7100
rect 35076 7044 35080 7100
rect 35016 7040 35080 7044
rect 35096 7100 35160 7104
rect 35096 7044 35100 7100
rect 35100 7044 35156 7100
rect 35156 7044 35160 7100
rect 35096 7040 35160 7044
rect 35176 7100 35240 7104
rect 35176 7044 35180 7100
rect 35180 7044 35236 7100
rect 35236 7044 35240 7100
rect 35176 7040 35240 7044
rect 19576 6556 19640 6560
rect 19576 6500 19580 6556
rect 19580 6500 19636 6556
rect 19636 6500 19640 6556
rect 19576 6496 19640 6500
rect 19656 6556 19720 6560
rect 19656 6500 19660 6556
rect 19660 6500 19716 6556
rect 19716 6500 19720 6556
rect 19656 6496 19720 6500
rect 19736 6556 19800 6560
rect 19736 6500 19740 6556
rect 19740 6500 19796 6556
rect 19796 6500 19800 6556
rect 19736 6496 19800 6500
rect 19816 6556 19880 6560
rect 19816 6500 19820 6556
rect 19820 6500 19876 6556
rect 19876 6500 19880 6556
rect 19816 6496 19880 6500
rect 50296 6556 50360 6560
rect 50296 6500 50300 6556
rect 50300 6500 50356 6556
rect 50356 6500 50360 6556
rect 50296 6496 50360 6500
rect 50376 6556 50440 6560
rect 50376 6500 50380 6556
rect 50380 6500 50436 6556
rect 50436 6500 50440 6556
rect 50376 6496 50440 6500
rect 50456 6556 50520 6560
rect 50456 6500 50460 6556
rect 50460 6500 50516 6556
rect 50516 6500 50520 6556
rect 50456 6496 50520 6500
rect 50536 6556 50600 6560
rect 50536 6500 50540 6556
rect 50540 6500 50596 6556
rect 50596 6500 50600 6556
rect 50536 6496 50600 6500
rect 4216 6012 4280 6016
rect 4216 5956 4220 6012
rect 4220 5956 4276 6012
rect 4276 5956 4280 6012
rect 4216 5952 4280 5956
rect 4296 6012 4360 6016
rect 4296 5956 4300 6012
rect 4300 5956 4356 6012
rect 4356 5956 4360 6012
rect 4296 5952 4360 5956
rect 4376 6012 4440 6016
rect 4376 5956 4380 6012
rect 4380 5956 4436 6012
rect 4436 5956 4440 6012
rect 4376 5952 4440 5956
rect 4456 6012 4520 6016
rect 4456 5956 4460 6012
rect 4460 5956 4516 6012
rect 4516 5956 4520 6012
rect 4456 5952 4520 5956
rect 34936 6012 35000 6016
rect 34936 5956 34940 6012
rect 34940 5956 34996 6012
rect 34996 5956 35000 6012
rect 34936 5952 35000 5956
rect 35016 6012 35080 6016
rect 35016 5956 35020 6012
rect 35020 5956 35076 6012
rect 35076 5956 35080 6012
rect 35016 5952 35080 5956
rect 35096 6012 35160 6016
rect 35096 5956 35100 6012
rect 35100 5956 35156 6012
rect 35156 5956 35160 6012
rect 35096 5952 35160 5956
rect 35176 6012 35240 6016
rect 35176 5956 35180 6012
rect 35180 5956 35236 6012
rect 35236 5956 35240 6012
rect 35176 5952 35240 5956
rect 19576 5468 19640 5472
rect 19576 5412 19580 5468
rect 19580 5412 19636 5468
rect 19636 5412 19640 5468
rect 19576 5408 19640 5412
rect 19656 5468 19720 5472
rect 19656 5412 19660 5468
rect 19660 5412 19716 5468
rect 19716 5412 19720 5468
rect 19656 5408 19720 5412
rect 19736 5468 19800 5472
rect 19736 5412 19740 5468
rect 19740 5412 19796 5468
rect 19796 5412 19800 5468
rect 19736 5408 19800 5412
rect 19816 5468 19880 5472
rect 19816 5412 19820 5468
rect 19820 5412 19876 5468
rect 19876 5412 19880 5468
rect 19816 5408 19880 5412
rect 50296 5468 50360 5472
rect 50296 5412 50300 5468
rect 50300 5412 50356 5468
rect 50356 5412 50360 5468
rect 50296 5408 50360 5412
rect 50376 5468 50440 5472
rect 50376 5412 50380 5468
rect 50380 5412 50436 5468
rect 50436 5412 50440 5468
rect 50376 5408 50440 5412
rect 50456 5468 50520 5472
rect 50456 5412 50460 5468
rect 50460 5412 50516 5468
rect 50516 5412 50520 5468
rect 50456 5408 50520 5412
rect 50536 5468 50600 5472
rect 50536 5412 50540 5468
rect 50540 5412 50596 5468
rect 50596 5412 50600 5468
rect 50536 5408 50600 5412
rect 4216 4924 4280 4928
rect 4216 4868 4220 4924
rect 4220 4868 4276 4924
rect 4276 4868 4280 4924
rect 4216 4864 4280 4868
rect 4296 4924 4360 4928
rect 4296 4868 4300 4924
rect 4300 4868 4356 4924
rect 4356 4868 4360 4924
rect 4296 4864 4360 4868
rect 4376 4924 4440 4928
rect 4376 4868 4380 4924
rect 4380 4868 4436 4924
rect 4436 4868 4440 4924
rect 4376 4864 4440 4868
rect 4456 4924 4520 4928
rect 4456 4868 4460 4924
rect 4460 4868 4516 4924
rect 4516 4868 4520 4924
rect 4456 4864 4520 4868
rect 34936 4924 35000 4928
rect 34936 4868 34940 4924
rect 34940 4868 34996 4924
rect 34996 4868 35000 4924
rect 34936 4864 35000 4868
rect 35016 4924 35080 4928
rect 35016 4868 35020 4924
rect 35020 4868 35076 4924
rect 35076 4868 35080 4924
rect 35016 4864 35080 4868
rect 35096 4924 35160 4928
rect 35096 4868 35100 4924
rect 35100 4868 35156 4924
rect 35156 4868 35160 4924
rect 35096 4864 35160 4868
rect 35176 4924 35240 4928
rect 35176 4868 35180 4924
rect 35180 4868 35236 4924
rect 35236 4868 35240 4924
rect 35176 4864 35240 4868
rect 19576 4380 19640 4384
rect 19576 4324 19580 4380
rect 19580 4324 19636 4380
rect 19636 4324 19640 4380
rect 19576 4320 19640 4324
rect 19656 4380 19720 4384
rect 19656 4324 19660 4380
rect 19660 4324 19716 4380
rect 19716 4324 19720 4380
rect 19656 4320 19720 4324
rect 19736 4380 19800 4384
rect 19736 4324 19740 4380
rect 19740 4324 19796 4380
rect 19796 4324 19800 4380
rect 19736 4320 19800 4324
rect 19816 4380 19880 4384
rect 19816 4324 19820 4380
rect 19820 4324 19876 4380
rect 19876 4324 19880 4380
rect 19816 4320 19880 4324
rect 50296 4380 50360 4384
rect 50296 4324 50300 4380
rect 50300 4324 50356 4380
rect 50356 4324 50360 4380
rect 50296 4320 50360 4324
rect 50376 4380 50440 4384
rect 50376 4324 50380 4380
rect 50380 4324 50436 4380
rect 50436 4324 50440 4380
rect 50376 4320 50440 4324
rect 50456 4380 50520 4384
rect 50456 4324 50460 4380
rect 50460 4324 50516 4380
rect 50516 4324 50520 4380
rect 50456 4320 50520 4324
rect 50536 4380 50600 4384
rect 50536 4324 50540 4380
rect 50540 4324 50596 4380
rect 50596 4324 50600 4380
rect 50536 4320 50600 4324
rect 4216 3836 4280 3840
rect 4216 3780 4220 3836
rect 4220 3780 4276 3836
rect 4276 3780 4280 3836
rect 4216 3776 4280 3780
rect 4296 3836 4360 3840
rect 4296 3780 4300 3836
rect 4300 3780 4356 3836
rect 4356 3780 4360 3836
rect 4296 3776 4360 3780
rect 4376 3836 4440 3840
rect 4376 3780 4380 3836
rect 4380 3780 4436 3836
rect 4436 3780 4440 3836
rect 4376 3776 4440 3780
rect 4456 3836 4520 3840
rect 4456 3780 4460 3836
rect 4460 3780 4516 3836
rect 4516 3780 4520 3836
rect 4456 3776 4520 3780
rect 34936 3836 35000 3840
rect 34936 3780 34940 3836
rect 34940 3780 34996 3836
rect 34996 3780 35000 3836
rect 34936 3776 35000 3780
rect 35016 3836 35080 3840
rect 35016 3780 35020 3836
rect 35020 3780 35076 3836
rect 35076 3780 35080 3836
rect 35016 3776 35080 3780
rect 35096 3836 35160 3840
rect 35096 3780 35100 3836
rect 35100 3780 35156 3836
rect 35156 3780 35160 3836
rect 35096 3776 35160 3780
rect 35176 3836 35240 3840
rect 35176 3780 35180 3836
rect 35180 3780 35236 3836
rect 35236 3780 35240 3836
rect 35176 3776 35240 3780
rect 19576 3292 19640 3296
rect 19576 3236 19580 3292
rect 19580 3236 19636 3292
rect 19636 3236 19640 3292
rect 19576 3232 19640 3236
rect 19656 3292 19720 3296
rect 19656 3236 19660 3292
rect 19660 3236 19716 3292
rect 19716 3236 19720 3292
rect 19656 3232 19720 3236
rect 19736 3292 19800 3296
rect 19736 3236 19740 3292
rect 19740 3236 19796 3292
rect 19796 3236 19800 3292
rect 19736 3232 19800 3236
rect 19816 3292 19880 3296
rect 19816 3236 19820 3292
rect 19820 3236 19876 3292
rect 19876 3236 19880 3292
rect 19816 3232 19880 3236
rect 50296 3292 50360 3296
rect 50296 3236 50300 3292
rect 50300 3236 50356 3292
rect 50356 3236 50360 3292
rect 50296 3232 50360 3236
rect 50376 3292 50440 3296
rect 50376 3236 50380 3292
rect 50380 3236 50436 3292
rect 50436 3236 50440 3292
rect 50376 3232 50440 3236
rect 50456 3292 50520 3296
rect 50456 3236 50460 3292
rect 50460 3236 50516 3292
rect 50516 3236 50520 3292
rect 50456 3232 50520 3236
rect 50536 3292 50600 3296
rect 50536 3236 50540 3292
rect 50540 3236 50596 3292
rect 50596 3236 50600 3292
rect 50536 3232 50600 3236
rect 4216 2748 4280 2752
rect 4216 2692 4220 2748
rect 4220 2692 4276 2748
rect 4276 2692 4280 2748
rect 4216 2688 4280 2692
rect 4296 2748 4360 2752
rect 4296 2692 4300 2748
rect 4300 2692 4356 2748
rect 4356 2692 4360 2748
rect 4296 2688 4360 2692
rect 4376 2748 4440 2752
rect 4376 2692 4380 2748
rect 4380 2692 4436 2748
rect 4436 2692 4440 2748
rect 4376 2688 4440 2692
rect 4456 2748 4520 2752
rect 4456 2692 4460 2748
rect 4460 2692 4516 2748
rect 4516 2692 4520 2748
rect 4456 2688 4520 2692
rect 34936 2748 35000 2752
rect 34936 2692 34940 2748
rect 34940 2692 34996 2748
rect 34996 2692 35000 2748
rect 34936 2688 35000 2692
rect 35016 2748 35080 2752
rect 35016 2692 35020 2748
rect 35020 2692 35076 2748
rect 35076 2692 35080 2748
rect 35016 2688 35080 2692
rect 35096 2748 35160 2752
rect 35096 2692 35100 2748
rect 35100 2692 35156 2748
rect 35156 2692 35160 2748
rect 35096 2688 35160 2692
rect 35176 2748 35240 2752
rect 35176 2692 35180 2748
rect 35180 2692 35236 2748
rect 35236 2692 35240 2748
rect 35176 2688 35240 2692
rect 19576 2204 19640 2208
rect 19576 2148 19580 2204
rect 19580 2148 19636 2204
rect 19636 2148 19640 2204
rect 19576 2144 19640 2148
rect 19656 2204 19720 2208
rect 19656 2148 19660 2204
rect 19660 2148 19716 2204
rect 19716 2148 19720 2204
rect 19656 2144 19720 2148
rect 19736 2204 19800 2208
rect 19736 2148 19740 2204
rect 19740 2148 19796 2204
rect 19796 2148 19800 2204
rect 19736 2144 19800 2148
rect 19816 2204 19880 2208
rect 19816 2148 19820 2204
rect 19820 2148 19876 2204
rect 19876 2148 19880 2204
rect 19816 2144 19880 2148
rect 50296 2204 50360 2208
rect 50296 2148 50300 2204
rect 50300 2148 50356 2204
rect 50356 2148 50360 2204
rect 50296 2144 50360 2148
rect 50376 2204 50440 2208
rect 50376 2148 50380 2204
rect 50380 2148 50436 2204
rect 50436 2148 50440 2204
rect 50376 2144 50440 2148
rect 50456 2204 50520 2208
rect 50456 2148 50460 2204
rect 50460 2148 50516 2204
rect 50516 2148 50520 2204
rect 50456 2144 50520 2148
rect 50536 2204 50600 2208
rect 50536 2148 50540 2204
rect 50540 2148 50596 2204
rect 50596 2148 50600 2204
rect 50536 2144 50600 2148
<< metal4 >>
rect 4208 57152 4528 57712
rect 4208 57088 4216 57152
rect 4280 57088 4296 57152
rect 4360 57088 4376 57152
rect 4440 57088 4456 57152
rect 4520 57088 4528 57152
rect 4208 56064 4528 57088
rect 4208 56000 4216 56064
rect 4280 56000 4296 56064
rect 4360 56000 4376 56064
rect 4440 56000 4456 56064
rect 4520 56000 4528 56064
rect 4208 54976 4528 56000
rect 4208 54912 4216 54976
rect 4280 54912 4296 54976
rect 4360 54912 4376 54976
rect 4440 54912 4456 54976
rect 4520 54912 4528 54976
rect 4208 53888 4528 54912
rect 4208 53824 4216 53888
rect 4280 53824 4296 53888
rect 4360 53824 4376 53888
rect 4440 53824 4456 53888
rect 4520 53824 4528 53888
rect 4208 52800 4528 53824
rect 4208 52736 4216 52800
rect 4280 52736 4296 52800
rect 4360 52736 4376 52800
rect 4440 52736 4456 52800
rect 4520 52736 4528 52800
rect 4208 51712 4528 52736
rect 4208 51648 4216 51712
rect 4280 51648 4296 51712
rect 4360 51648 4376 51712
rect 4440 51648 4456 51712
rect 4520 51648 4528 51712
rect 4208 50624 4528 51648
rect 4208 50560 4216 50624
rect 4280 50560 4296 50624
rect 4360 50560 4376 50624
rect 4440 50560 4456 50624
rect 4520 50560 4528 50624
rect 4208 49536 4528 50560
rect 4208 49472 4216 49536
rect 4280 49472 4296 49536
rect 4360 49472 4376 49536
rect 4440 49472 4456 49536
rect 4520 49472 4528 49536
rect 4208 48448 4528 49472
rect 4208 48384 4216 48448
rect 4280 48384 4296 48448
rect 4360 48384 4376 48448
rect 4440 48384 4456 48448
rect 4520 48384 4528 48448
rect 4208 47360 4528 48384
rect 4208 47296 4216 47360
rect 4280 47296 4296 47360
rect 4360 47296 4376 47360
rect 4440 47296 4456 47360
rect 4520 47296 4528 47360
rect 4208 46272 4528 47296
rect 4208 46208 4216 46272
rect 4280 46208 4296 46272
rect 4360 46208 4376 46272
rect 4440 46208 4456 46272
rect 4520 46208 4528 46272
rect 4208 45184 4528 46208
rect 4208 45120 4216 45184
rect 4280 45120 4296 45184
rect 4360 45120 4376 45184
rect 4440 45120 4456 45184
rect 4520 45120 4528 45184
rect 4208 44096 4528 45120
rect 4208 44032 4216 44096
rect 4280 44032 4296 44096
rect 4360 44032 4376 44096
rect 4440 44032 4456 44096
rect 4520 44032 4528 44096
rect 4208 43008 4528 44032
rect 4208 42944 4216 43008
rect 4280 42944 4296 43008
rect 4360 42944 4376 43008
rect 4440 42944 4456 43008
rect 4520 42944 4528 43008
rect 4208 41920 4528 42944
rect 4208 41856 4216 41920
rect 4280 41856 4296 41920
rect 4360 41856 4376 41920
rect 4440 41856 4456 41920
rect 4520 41856 4528 41920
rect 4208 40832 4528 41856
rect 4208 40768 4216 40832
rect 4280 40768 4296 40832
rect 4360 40768 4376 40832
rect 4440 40768 4456 40832
rect 4520 40768 4528 40832
rect 4208 39744 4528 40768
rect 4208 39680 4216 39744
rect 4280 39680 4296 39744
rect 4360 39680 4376 39744
rect 4440 39680 4456 39744
rect 4520 39680 4528 39744
rect 4208 38656 4528 39680
rect 4208 38592 4216 38656
rect 4280 38592 4296 38656
rect 4360 38592 4376 38656
rect 4440 38592 4456 38656
rect 4520 38592 4528 38656
rect 4208 37568 4528 38592
rect 4208 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4528 37568
rect 4208 36480 4528 37504
rect 4208 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4528 36480
rect 4208 35392 4528 36416
rect 4208 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4528 35392
rect 4208 34304 4528 35328
rect 4208 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4528 34304
rect 4208 33216 4528 34240
rect 4208 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4528 33216
rect 4208 32128 4528 33152
rect 4208 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4528 32128
rect 4208 31040 4528 32064
rect 4208 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4528 31040
rect 4208 29952 4528 30976
rect 4208 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4528 29952
rect 4208 28864 4528 29888
rect 4208 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4528 28864
rect 4208 27776 4528 28800
rect 4208 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4528 27776
rect 4208 26688 4528 27712
rect 4208 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4528 26688
rect 4208 25600 4528 26624
rect 4208 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4528 25600
rect 4208 24512 4528 25536
rect 4208 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4528 24512
rect 4208 23424 4528 24448
rect 4208 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4528 23424
rect 4208 22336 4528 23360
rect 4208 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4528 22336
rect 4208 21248 4528 22272
rect 4208 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4528 21248
rect 4208 20160 4528 21184
rect 4208 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4528 20160
rect 4208 19072 4528 20096
rect 4208 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4528 19072
rect 4208 17984 4528 19008
rect 4208 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4528 17984
rect 4208 16896 4528 17920
rect 4208 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4528 16896
rect 4208 15808 4528 16832
rect 4208 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4528 15808
rect 4208 14720 4528 15744
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 4208 13632 4528 14656
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 12544 4528 13568
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 11456 4528 12480
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 10368 4528 11392
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 9280 4528 10304
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 8192 4528 9216
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 7104 4528 8128
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 6016 4528 7040
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 4928 4528 5952
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 3840 4528 4864
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 2752 4528 3776
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2128 4528 2688
rect 19568 57696 19888 57712
rect 19568 57632 19576 57696
rect 19640 57632 19656 57696
rect 19720 57632 19736 57696
rect 19800 57632 19816 57696
rect 19880 57632 19888 57696
rect 19568 56608 19888 57632
rect 19568 56544 19576 56608
rect 19640 56544 19656 56608
rect 19720 56544 19736 56608
rect 19800 56544 19816 56608
rect 19880 56544 19888 56608
rect 19568 55520 19888 56544
rect 19568 55456 19576 55520
rect 19640 55456 19656 55520
rect 19720 55456 19736 55520
rect 19800 55456 19816 55520
rect 19880 55456 19888 55520
rect 19568 54432 19888 55456
rect 19568 54368 19576 54432
rect 19640 54368 19656 54432
rect 19720 54368 19736 54432
rect 19800 54368 19816 54432
rect 19880 54368 19888 54432
rect 19568 53344 19888 54368
rect 19568 53280 19576 53344
rect 19640 53280 19656 53344
rect 19720 53280 19736 53344
rect 19800 53280 19816 53344
rect 19880 53280 19888 53344
rect 19568 52256 19888 53280
rect 19568 52192 19576 52256
rect 19640 52192 19656 52256
rect 19720 52192 19736 52256
rect 19800 52192 19816 52256
rect 19880 52192 19888 52256
rect 19568 51168 19888 52192
rect 19568 51104 19576 51168
rect 19640 51104 19656 51168
rect 19720 51104 19736 51168
rect 19800 51104 19816 51168
rect 19880 51104 19888 51168
rect 19568 50080 19888 51104
rect 19568 50016 19576 50080
rect 19640 50016 19656 50080
rect 19720 50016 19736 50080
rect 19800 50016 19816 50080
rect 19880 50016 19888 50080
rect 19568 48992 19888 50016
rect 19568 48928 19576 48992
rect 19640 48928 19656 48992
rect 19720 48928 19736 48992
rect 19800 48928 19816 48992
rect 19880 48928 19888 48992
rect 19568 47904 19888 48928
rect 19568 47840 19576 47904
rect 19640 47840 19656 47904
rect 19720 47840 19736 47904
rect 19800 47840 19816 47904
rect 19880 47840 19888 47904
rect 19568 46816 19888 47840
rect 19568 46752 19576 46816
rect 19640 46752 19656 46816
rect 19720 46752 19736 46816
rect 19800 46752 19816 46816
rect 19880 46752 19888 46816
rect 19568 45728 19888 46752
rect 19568 45664 19576 45728
rect 19640 45664 19656 45728
rect 19720 45664 19736 45728
rect 19800 45664 19816 45728
rect 19880 45664 19888 45728
rect 19568 44640 19888 45664
rect 19568 44576 19576 44640
rect 19640 44576 19656 44640
rect 19720 44576 19736 44640
rect 19800 44576 19816 44640
rect 19880 44576 19888 44640
rect 19568 43552 19888 44576
rect 19568 43488 19576 43552
rect 19640 43488 19656 43552
rect 19720 43488 19736 43552
rect 19800 43488 19816 43552
rect 19880 43488 19888 43552
rect 19568 42464 19888 43488
rect 19568 42400 19576 42464
rect 19640 42400 19656 42464
rect 19720 42400 19736 42464
rect 19800 42400 19816 42464
rect 19880 42400 19888 42464
rect 19568 41376 19888 42400
rect 19568 41312 19576 41376
rect 19640 41312 19656 41376
rect 19720 41312 19736 41376
rect 19800 41312 19816 41376
rect 19880 41312 19888 41376
rect 19568 40288 19888 41312
rect 19568 40224 19576 40288
rect 19640 40224 19656 40288
rect 19720 40224 19736 40288
rect 19800 40224 19816 40288
rect 19880 40224 19888 40288
rect 19568 39200 19888 40224
rect 19568 39136 19576 39200
rect 19640 39136 19656 39200
rect 19720 39136 19736 39200
rect 19800 39136 19816 39200
rect 19880 39136 19888 39200
rect 19568 38112 19888 39136
rect 19568 38048 19576 38112
rect 19640 38048 19656 38112
rect 19720 38048 19736 38112
rect 19800 38048 19816 38112
rect 19880 38048 19888 38112
rect 19568 37024 19888 38048
rect 19568 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19888 37024
rect 19568 35936 19888 36960
rect 19568 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19888 35936
rect 19568 34848 19888 35872
rect 19568 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19888 34848
rect 19568 33760 19888 34784
rect 19568 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19888 33760
rect 19568 32672 19888 33696
rect 19568 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19888 32672
rect 19568 31584 19888 32608
rect 19568 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19888 31584
rect 19568 30496 19888 31520
rect 19568 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19888 30496
rect 19568 29408 19888 30432
rect 19568 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19888 29408
rect 19568 28320 19888 29344
rect 19568 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19888 28320
rect 19568 27232 19888 28256
rect 19568 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19888 27232
rect 19568 26144 19888 27168
rect 19568 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19888 26144
rect 19568 25056 19888 26080
rect 19568 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19888 25056
rect 19568 23968 19888 24992
rect 19568 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19888 23968
rect 19568 22880 19888 23904
rect 19568 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19888 22880
rect 19568 21792 19888 22816
rect 19568 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19888 21792
rect 19568 20704 19888 21728
rect 19568 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19888 20704
rect 19568 19616 19888 20640
rect 19568 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19888 19616
rect 19568 18528 19888 19552
rect 19568 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19888 18528
rect 19568 17440 19888 18464
rect 19568 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19888 17440
rect 19568 16352 19888 17376
rect 19568 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19888 16352
rect 19568 15264 19888 16288
rect 19568 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19888 15264
rect 19568 14176 19888 15200
rect 19568 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19888 14176
rect 19568 13088 19888 14112
rect 19568 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19888 13088
rect 19568 12000 19888 13024
rect 19568 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19888 12000
rect 19568 10912 19888 11936
rect 19568 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19888 10912
rect 19568 9824 19888 10848
rect 19568 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19888 9824
rect 19568 8736 19888 9760
rect 19568 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19888 8736
rect 19568 7648 19888 8672
rect 19568 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19888 7648
rect 19568 6560 19888 7584
rect 19568 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19888 6560
rect 19568 5472 19888 6496
rect 19568 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19888 5472
rect 19568 4384 19888 5408
rect 19568 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19888 4384
rect 19568 3296 19888 4320
rect 19568 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19888 3296
rect 19568 2208 19888 3232
rect 19568 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19888 2208
rect 19568 2128 19888 2144
rect 34928 57152 35248 57712
rect 34928 57088 34936 57152
rect 35000 57088 35016 57152
rect 35080 57088 35096 57152
rect 35160 57088 35176 57152
rect 35240 57088 35248 57152
rect 34928 56064 35248 57088
rect 34928 56000 34936 56064
rect 35000 56000 35016 56064
rect 35080 56000 35096 56064
rect 35160 56000 35176 56064
rect 35240 56000 35248 56064
rect 34928 54976 35248 56000
rect 34928 54912 34936 54976
rect 35000 54912 35016 54976
rect 35080 54912 35096 54976
rect 35160 54912 35176 54976
rect 35240 54912 35248 54976
rect 34928 53888 35248 54912
rect 34928 53824 34936 53888
rect 35000 53824 35016 53888
rect 35080 53824 35096 53888
rect 35160 53824 35176 53888
rect 35240 53824 35248 53888
rect 34928 52800 35248 53824
rect 34928 52736 34936 52800
rect 35000 52736 35016 52800
rect 35080 52736 35096 52800
rect 35160 52736 35176 52800
rect 35240 52736 35248 52800
rect 34928 51712 35248 52736
rect 34928 51648 34936 51712
rect 35000 51648 35016 51712
rect 35080 51648 35096 51712
rect 35160 51648 35176 51712
rect 35240 51648 35248 51712
rect 34928 50624 35248 51648
rect 34928 50560 34936 50624
rect 35000 50560 35016 50624
rect 35080 50560 35096 50624
rect 35160 50560 35176 50624
rect 35240 50560 35248 50624
rect 34928 49536 35248 50560
rect 34928 49472 34936 49536
rect 35000 49472 35016 49536
rect 35080 49472 35096 49536
rect 35160 49472 35176 49536
rect 35240 49472 35248 49536
rect 34928 48448 35248 49472
rect 34928 48384 34936 48448
rect 35000 48384 35016 48448
rect 35080 48384 35096 48448
rect 35160 48384 35176 48448
rect 35240 48384 35248 48448
rect 34928 47360 35248 48384
rect 34928 47296 34936 47360
rect 35000 47296 35016 47360
rect 35080 47296 35096 47360
rect 35160 47296 35176 47360
rect 35240 47296 35248 47360
rect 34928 46272 35248 47296
rect 34928 46208 34936 46272
rect 35000 46208 35016 46272
rect 35080 46208 35096 46272
rect 35160 46208 35176 46272
rect 35240 46208 35248 46272
rect 34928 45184 35248 46208
rect 34928 45120 34936 45184
rect 35000 45120 35016 45184
rect 35080 45120 35096 45184
rect 35160 45120 35176 45184
rect 35240 45120 35248 45184
rect 34928 44096 35248 45120
rect 34928 44032 34936 44096
rect 35000 44032 35016 44096
rect 35080 44032 35096 44096
rect 35160 44032 35176 44096
rect 35240 44032 35248 44096
rect 34928 43008 35248 44032
rect 34928 42944 34936 43008
rect 35000 42944 35016 43008
rect 35080 42944 35096 43008
rect 35160 42944 35176 43008
rect 35240 42944 35248 43008
rect 34928 41920 35248 42944
rect 34928 41856 34936 41920
rect 35000 41856 35016 41920
rect 35080 41856 35096 41920
rect 35160 41856 35176 41920
rect 35240 41856 35248 41920
rect 34928 40832 35248 41856
rect 34928 40768 34936 40832
rect 35000 40768 35016 40832
rect 35080 40768 35096 40832
rect 35160 40768 35176 40832
rect 35240 40768 35248 40832
rect 34928 39744 35248 40768
rect 34928 39680 34936 39744
rect 35000 39680 35016 39744
rect 35080 39680 35096 39744
rect 35160 39680 35176 39744
rect 35240 39680 35248 39744
rect 34928 38656 35248 39680
rect 34928 38592 34936 38656
rect 35000 38592 35016 38656
rect 35080 38592 35096 38656
rect 35160 38592 35176 38656
rect 35240 38592 35248 38656
rect 34928 37568 35248 38592
rect 34928 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35248 37568
rect 34928 36480 35248 37504
rect 34928 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35248 36480
rect 34928 35392 35248 36416
rect 34928 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35248 35392
rect 34928 34304 35248 35328
rect 34928 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35248 34304
rect 34928 33216 35248 34240
rect 34928 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35248 33216
rect 34928 32128 35248 33152
rect 34928 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35248 32128
rect 34928 31040 35248 32064
rect 34928 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35248 31040
rect 34928 29952 35248 30976
rect 34928 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35248 29952
rect 34928 28864 35248 29888
rect 34928 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35248 28864
rect 34928 27776 35248 28800
rect 34928 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35248 27776
rect 34928 26688 35248 27712
rect 34928 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35248 26688
rect 34928 25600 35248 26624
rect 34928 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35248 25600
rect 34928 24512 35248 25536
rect 34928 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35248 24512
rect 34928 23424 35248 24448
rect 34928 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35248 23424
rect 34928 22336 35248 23360
rect 34928 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35248 22336
rect 34928 21248 35248 22272
rect 34928 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35248 21248
rect 34928 20160 35248 21184
rect 34928 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35248 20160
rect 34928 19072 35248 20096
rect 34928 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35248 19072
rect 34928 17984 35248 19008
rect 34928 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35248 17984
rect 34928 16896 35248 17920
rect 34928 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35248 16896
rect 34928 15808 35248 16832
rect 34928 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35248 15808
rect 34928 14720 35248 15744
rect 34928 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35248 14720
rect 34928 13632 35248 14656
rect 34928 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35248 13632
rect 34928 12544 35248 13568
rect 34928 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35248 12544
rect 34928 11456 35248 12480
rect 34928 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35248 11456
rect 34928 10368 35248 11392
rect 34928 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35248 10368
rect 34928 9280 35248 10304
rect 34928 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35248 9280
rect 34928 8192 35248 9216
rect 34928 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35248 8192
rect 34928 7104 35248 8128
rect 34928 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35248 7104
rect 34928 6016 35248 7040
rect 34928 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35248 6016
rect 34928 4928 35248 5952
rect 34928 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35248 4928
rect 34928 3840 35248 4864
rect 34928 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35248 3840
rect 34928 2752 35248 3776
rect 34928 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35248 2752
rect 34928 2128 35248 2688
rect 50288 57696 50608 57712
rect 50288 57632 50296 57696
rect 50360 57632 50376 57696
rect 50440 57632 50456 57696
rect 50520 57632 50536 57696
rect 50600 57632 50608 57696
rect 50288 56608 50608 57632
rect 50288 56544 50296 56608
rect 50360 56544 50376 56608
rect 50440 56544 50456 56608
rect 50520 56544 50536 56608
rect 50600 56544 50608 56608
rect 50288 55520 50608 56544
rect 50288 55456 50296 55520
rect 50360 55456 50376 55520
rect 50440 55456 50456 55520
rect 50520 55456 50536 55520
rect 50600 55456 50608 55520
rect 50288 54432 50608 55456
rect 50288 54368 50296 54432
rect 50360 54368 50376 54432
rect 50440 54368 50456 54432
rect 50520 54368 50536 54432
rect 50600 54368 50608 54432
rect 50288 53344 50608 54368
rect 50288 53280 50296 53344
rect 50360 53280 50376 53344
rect 50440 53280 50456 53344
rect 50520 53280 50536 53344
rect 50600 53280 50608 53344
rect 50288 52256 50608 53280
rect 50288 52192 50296 52256
rect 50360 52192 50376 52256
rect 50440 52192 50456 52256
rect 50520 52192 50536 52256
rect 50600 52192 50608 52256
rect 50288 51168 50608 52192
rect 50288 51104 50296 51168
rect 50360 51104 50376 51168
rect 50440 51104 50456 51168
rect 50520 51104 50536 51168
rect 50600 51104 50608 51168
rect 50288 50080 50608 51104
rect 50288 50016 50296 50080
rect 50360 50016 50376 50080
rect 50440 50016 50456 50080
rect 50520 50016 50536 50080
rect 50600 50016 50608 50080
rect 50288 48992 50608 50016
rect 50288 48928 50296 48992
rect 50360 48928 50376 48992
rect 50440 48928 50456 48992
rect 50520 48928 50536 48992
rect 50600 48928 50608 48992
rect 50288 47904 50608 48928
rect 50288 47840 50296 47904
rect 50360 47840 50376 47904
rect 50440 47840 50456 47904
rect 50520 47840 50536 47904
rect 50600 47840 50608 47904
rect 50288 46816 50608 47840
rect 50288 46752 50296 46816
rect 50360 46752 50376 46816
rect 50440 46752 50456 46816
rect 50520 46752 50536 46816
rect 50600 46752 50608 46816
rect 50288 45728 50608 46752
rect 50288 45664 50296 45728
rect 50360 45664 50376 45728
rect 50440 45664 50456 45728
rect 50520 45664 50536 45728
rect 50600 45664 50608 45728
rect 50288 44640 50608 45664
rect 50288 44576 50296 44640
rect 50360 44576 50376 44640
rect 50440 44576 50456 44640
rect 50520 44576 50536 44640
rect 50600 44576 50608 44640
rect 50288 43552 50608 44576
rect 50288 43488 50296 43552
rect 50360 43488 50376 43552
rect 50440 43488 50456 43552
rect 50520 43488 50536 43552
rect 50600 43488 50608 43552
rect 50288 42464 50608 43488
rect 50288 42400 50296 42464
rect 50360 42400 50376 42464
rect 50440 42400 50456 42464
rect 50520 42400 50536 42464
rect 50600 42400 50608 42464
rect 50288 41376 50608 42400
rect 50288 41312 50296 41376
rect 50360 41312 50376 41376
rect 50440 41312 50456 41376
rect 50520 41312 50536 41376
rect 50600 41312 50608 41376
rect 50288 40288 50608 41312
rect 50288 40224 50296 40288
rect 50360 40224 50376 40288
rect 50440 40224 50456 40288
rect 50520 40224 50536 40288
rect 50600 40224 50608 40288
rect 50288 39200 50608 40224
rect 50288 39136 50296 39200
rect 50360 39136 50376 39200
rect 50440 39136 50456 39200
rect 50520 39136 50536 39200
rect 50600 39136 50608 39200
rect 50288 38112 50608 39136
rect 50288 38048 50296 38112
rect 50360 38048 50376 38112
rect 50440 38048 50456 38112
rect 50520 38048 50536 38112
rect 50600 38048 50608 38112
rect 50288 37024 50608 38048
rect 50288 36960 50296 37024
rect 50360 36960 50376 37024
rect 50440 36960 50456 37024
rect 50520 36960 50536 37024
rect 50600 36960 50608 37024
rect 50288 35936 50608 36960
rect 50288 35872 50296 35936
rect 50360 35872 50376 35936
rect 50440 35872 50456 35936
rect 50520 35872 50536 35936
rect 50600 35872 50608 35936
rect 50288 34848 50608 35872
rect 50288 34784 50296 34848
rect 50360 34784 50376 34848
rect 50440 34784 50456 34848
rect 50520 34784 50536 34848
rect 50600 34784 50608 34848
rect 50288 33760 50608 34784
rect 50288 33696 50296 33760
rect 50360 33696 50376 33760
rect 50440 33696 50456 33760
rect 50520 33696 50536 33760
rect 50600 33696 50608 33760
rect 50288 32672 50608 33696
rect 50288 32608 50296 32672
rect 50360 32608 50376 32672
rect 50440 32608 50456 32672
rect 50520 32608 50536 32672
rect 50600 32608 50608 32672
rect 50288 31584 50608 32608
rect 50288 31520 50296 31584
rect 50360 31520 50376 31584
rect 50440 31520 50456 31584
rect 50520 31520 50536 31584
rect 50600 31520 50608 31584
rect 50288 30496 50608 31520
rect 50288 30432 50296 30496
rect 50360 30432 50376 30496
rect 50440 30432 50456 30496
rect 50520 30432 50536 30496
rect 50600 30432 50608 30496
rect 50288 29408 50608 30432
rect 50288 29344 50296 29408
rect 50360 29344 50376 29408
rect 50440 29344 50456 29408
rect 50520 29344 50536 29408
rect 50600 29344 50608 29408
rect 50288 28320 50608 29344
rect 50288 28256 50296 28320
rect 50360 28256 50376 28320
rect 50440 28256 50456 28320
rect 50520 28256 50536 28320
rect 50600 28256 50608 28320
rect 50288 27232 50608 28256
rect 50288 27168 50296 27232
rect 50360 27168 50376 27232
rect 50440 27168 50456 27232
rect 50520 27168 50536 27232
rect 50600 27168 50608 27232
rect 50288 26144 50608 27168
rect 50288 26080 50296 26144
rect 50360 26080 50376 26144
rect 50440 26080 50456 26144
rect 50520 26080 50536 26144
rect 50600 26080 50608 26144
rect 50288 25056 50608 26080
rect 50288 24992 50296 25056
rect 50360 24992 50376 25056
rect 50440 24992 50456 25056
rect 50520 24992 50536 25056
rect 50600 24992 50608 25056
rect 50288 23968 50608 24992
rect 50288 23904 50296 23968
rect 50360 23904 50376 23968
rect 50440 23904 50456 23968
rect 50520 23904 50536 23968
rect 50600 23904 50608 23968
rect 50288 22880 50608 23904
rect 50288 22816 50296 22880
rect 50360 22816 50376 22880
rect 50440 22816 50456 22880
rect 50520 22816 50536 22880
rect 50600 22816 50608 22880
rect 50288 21792 50608 22816
rect 50288 21728 50296 21792
rect 50360 21728 50376 21792
rect 50440 21728 50456 21792
rect 50520 21728 50536 21792
rect 50600 21728 50608 21792
rect 50288 20704 50608 21728
rect 50288 20640 50296 20704
rect 50360 20640 50376 20704
rect 50440 20640 50456 20704
rect 50520 20640 50536 20704
rect 50600 20640 50608 20704
rect 50288 19616 50608 20640
rect 50288 19552 50296 19616
rect 50360 19552 50376 19616
rect 50440 19552 50456 19616
rect 50520 19552 50536 19616
rect 50600 19552 50608 19616
rect 50288 18528 50608 19552
rect 50288 18464 50296 18528
rect 50360 18464 50376 18528
rect 50440 18464 50456 18528
rect 50520 18464 50536 18528
rect 50600 18464 50608 18528
rect 50288 17440 50608 18464
rect 50288 17376 50296 17440
rect 50360 17376 50376 17440
rect 50440 17376 50456 17440
rect 50520 17376 50536 17440
rect 50600 17376 50608 17440
rect 50288 16352 50608 17376
rect 50288 16288 50296 16352
rect 50360 16288 50376 16352
rect 50440 16288 50456 16352
rect 50520 16288 50536 16352
rect 50600 16288 50608 16352
rect 50288 15264 50608 16288
rect 50288 15200 50296 15264
rect 50360 15200 50376 15264
rect 50440 15200 50456 15264
rect 50520 15200 50536 15264
rect 50600 15200 50608 15264
rect 50288 14176 50608 15200
rect 50288 14112 50296 14176
rect 50360 14112 50376 14176
rect 50440 14112 50456 14176
rect 50520 14112 50536 14176
rect 50600 14112 50608 14176
rect 50288 13088 50608 14112
rect 50288 13024 50296 13088
rect 50360 13024 50376 13088
rect 50440 13024 50456 13088
rect 50520 13024 50536 13088
rect 50600 13024 50608 13088
rect 50288 12000 50608 13024
rect 50288 11936 50296 12000
rect 50360 11936 50376 12000
rect 50440 11936 50456 12000
rect 50520 11936 50536 12000
rect 50600 11936 50608 12000
rect 50288 10912 50608 11936
rect 50288 10848 50296 10912
rect 50360 10848 50376 10912
rect 50440 10848 50456 10912
rect 50520 10848 50536 10912
rect 50600 10848 50608 10912
rect 50288 9824 50608 10848
rect 50288 9760 50296 9824
rect 50360 9760 50376 9824
rect 50440 9760 50456 9824
rect 50520 9760 50536 9824
rect 50600 9760 50608 9824
rect 50288 8736 50608 9760
rect 50288 8672 50296 8736
rect 50360 8672 50376 8736
rect 50440 8672 50456 8736
rect 50520 8672 50536 8736
rect 50600 8672 50608 8736
rect 50288 7648 50608 8672
rect 50288 7584 50296 7648
rect 50360 7584 50376 7648
rect 50440 7584 50456 7648
rect 50520 7584 50536 7648
rect 50600 7584 50608 7648
rect 50288 6560 50608 7584
rect 50288 6496 50296 6560
rect 50360 6496 50376 6560
rect 50440 6496 50456 6560
rect 50520 6496 50536 6560
rect 50600 6496 50608 6560
rect 50288 5472 50608 6496
rect 50288 5408 50296 5472
rect 50360 5408 50376 5472
rect 50440 5408 50456 5472
rect 50520 5408 50536 5472
rect 50600 5408 50608 5472
rect 50288 4384 50608 5408
rect 50288 4320 50296 4384
rect 50360 4320 50376 4384
rect 50440 4320 50456 4384
rect 50520 4320 50536 4384
rect 50600 4320 50608 4384
rect 50288 3296 50608 4320
rect 50288 3232 50296 3296
rect 50360 3232 50376 3296
rect 50440 3232 50456 3296
rect 50520 3232 50536 3296
rect 50600 3232 50608 3296
rect 50288 2208 50608 3232
rect 50288 2144 50296 2208
rect 50360 2144 50376 2208
rect 50440 2144 50456 2208
rect 50520 2144 50536 2208
rect 50600 2144 50608 2208
rect 50288 2128 50608 2144
use sky130_fd_sc_hd__decap_12  FILLER_0_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 1380 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_15
timestamp 1644511149
transform 1 0 2484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_29
timestamp 1644511149
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_41
timestamp 1644511149
transform 1 0 4876 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 5980 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_57 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 6348 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_65
timestamp 1644511149
transform 1 0 7084 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_72
timestamp 1644511149
transform 1 0 7728 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_85
timestamp 1644511149
transform 1 0 8924 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_97
timestamp 1644511149
transform 1 0 10028 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_109
timestamp 1644511149
transform 1 0 11132 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_113
timestamp 1644511149
transform 1 0 11500 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_125
timestamp 1644511149
transform 1 0 12604 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_137
timestamp 1644511149
transform 1 0 13708 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_141
timestamp 1644511149
transform 1 0 14076 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_153
timestamp 1644511149
transform 1 0 15180 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_165
timestamp 1644511149
transform 1 0 16284 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_169
timestamp 1644511149
transform 1 0 16652 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_181
timestamp 1644511149
transform 1 0 17756 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_193
timestamp 1644511149
transform 1 0 18860 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_197
timestamp 1644511149
transform 1 0 19228 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_209
timestamp 1644511149
transform 1 0 20332 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_221
timestamp 1644511149
transform 1 0 21436 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_225
timestamp 1644511149
transform 1 0 21804 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_237
timestamp 1644511149
transform 1 0 22908 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_249
timestamp 1644511149
transform 1 0 24012 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_262
timestamp 1644511149
transform 1 0 25208 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_274 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 26312 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_281
timestamp 1644511149
transform 1 0 26956 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_293
timestamp 1644511149
transform 1 0 28060 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_305
timestamp 1644511149
transform 1 0 29164 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_309
timestamp 1644511149
transform 1 0 29532 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_321
timestamp 1644511149
transform 1 0 30636 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_333
timestamp 1644511149
transform 1 0 31740 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_337
timestamp 1644511149
transform 1 0 32108 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_349
timestamp 1644511149
transform 1 0 33212 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_361
timestamp 1644511149
transform 1 0 34316 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_365
timestamp 1644511149
transform 1 0 34684 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_377
timestamp 1644511149
transform 1 0 35788 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_389
timestamp 1644511149
transform 1 0 36892 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_393
timestamp 1644511149
transform 1 0 37260 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_405
timestamp 1644511149
transform 1 0 38364 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_417
timestamp 1644511149
transform 1 0 39468 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_421
timestamp 1644511149
transform 1 0 39836 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_433
timestamp 1644511149
transform 1 0 40940 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_445
timestamp 1644511149
transform 1 0 42044 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_449
timestamp 1644511149
transform 1 0 42412 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_461
timestamp 1644511149
transform 1 0 43516 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_473
timestamp 1644511149
transform 1 0 44620 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_477
timestamp 1644511149
transform 1 0 44988 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_489
timestamp 1644511149
transform 1 0 46092 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_501
timestamp 1644511149
transform 1 0 47196 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_505
timestamp 1644511149
transform 1 0 47564 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_517
timestamp 1644511149
transform 1 0 48668 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_529
timestamp 1644511149
transform 1 0 49772 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_533
timestamp 1644511149
transform 1 0 50140 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_545
timestamp 1644511149
transform 1 0 51244 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_557
timestamp 1644511149
transform 1 0 52348 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_561
timestamp 1644511149
transform 1 0 52716 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_573
timestamp 1644511149
transform 1 0 53820 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_585
timestamp 1644511149
transform 1 0 54924 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_589
timestamp 1644511149
transform 1 0 55292 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_601 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 56396 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_606
timestamp 1644511149
transform 1 0 56856 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_614
timestamp 1644511149
transform 1 0 57592 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_620 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 58144 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_624
timestamp 1644511149
transform 1 0 58512 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_3
timestamp 1644511149
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_15
timestamp 1644511149
transform 1 0 2484 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_27
timestamp 1644511149
transform 1 0 3588 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_1_36
timestamp 1644511149
transform 1 0 4416 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_48
timestamp 1644511149
transform 1 0 5520 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_1_57
timestamp 1644511149
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_69
timestamp 1644511149
transform 1 0 7452 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_81
timestamp 1644511149
transform 1 0 8556 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_93
timestamp 1644511149
transform 1 0 9660 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_105
timestamp 1644511149
transform 1 0 10764 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_111
timestamp 1644511149
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_113
timestamp 1644511149
transform 1 0 11500 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_125
timestamp 1644511149
transform 1 0 12604 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_137
timestamp 1644511149
transform 1 0 13708 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_1_148
timestamp 1644511149
transform 1 0 14720 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_154
timestamp 1644511149
transform 1 0 15272 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_158
timestamp 1644511149
transform 1 0 15640 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_166
timestamp 1644511149
transform 1 0 16376 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_1_169
timestamp 1644511149
transform 1 0 16652 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_1_178
timestamp 1644511149
transform 1 0 17480 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_186
timestamp 1644511149
transform 1 0 18216 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_190
timestamp 1644511149
transform 1 0 18584 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_202
timestamp 1644511149
transform 1 0 19688 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_1_210
timestamp 1644511149
transform 1 0 20424 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_1_216
timestamp 1644511149
transform 1 0 20976 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_1_225
timestamp 1644511149
transform 1 0 21804 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_237
timestamp 1644511149
transform 1 0 22908 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_249
timestamp 1644511149
transform 1 0 24012 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_261
timestamp 1644511149
transform 1 0 25116 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_273
timestamp 1644511149
transform 1 0 26220 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_279
timestamp 1644511149
transform 1 0 26772 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_281
timestamp 1644511149
transform 1 0 26956 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_293
timestamp 1644511149
transform 1 0 28060 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_305
timestamp 1644511149
transform 1 0 29164 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_317
timestamp 1644511149
transform 1 0 30268 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_329
timestamp 1644511149
transform 1 0 31372 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_335
timestamp 1644511149
transform 1 0 31924 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_337
timestamp 1644511149
transform 1 0 32108 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_349
timestamp 1644511149
transform 1 0 33212 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_361
timestamp 1644511149
transform 1 0 34316 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_373
timestamp 1644511149
transform 1 0 35420 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_385
timestamp 1644511149
transform 1 0 36524 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_391
timestamp 1644511149
transform 1 0 37076 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_393
timestamp 1644511149
transform 1 0 37260 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_405
timestamp 1644511149
transform 1 0 38364 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_417
timestamp 1644511149
transform 1 0 39468 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_429
timestamp 1644511149
transform 1 0 40572 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_441
timestamp 1644511149
transform 1 0 41676 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_447
timestamp 1644511149
transform 1 0 42228 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_449
timestamp 1644511149
transform 1 0 42412 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_461
timestamp 1644511149
transform 1 0 43516 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_469
timestamp 1644511149
transform 1 0 44252 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_1_474
timestamp 1644511149
transform 1 0 44712 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_486
timestamp 1644511149
transform 1 0 45816 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_498
timestamp 1644511149
transform 1 0 46920 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_1_505
timestamp 1644511149
transform 1 0 47564 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_517
timestamp 1644511149
transform 1 0 48668 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_529
timestamp 1644511149
transform 1 0 49772 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_541
timestamp 1644511149
transform 1 0 50876 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_547
timestamp 1644511149
transform 1 0 51428 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_551
timestamp 1644511149
transform 1 0 51796 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_559
timestamp 1644511149
transform 1 0 52532 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_561
timestamp 1644511149
transform 1 0 52716 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_573
timestamp 1644511149
transform 1 0 53820 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_579
timestamp 1644511149
transform 1 0 54372 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_601
timestamp 1644511149
transform 1 0 56396 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_608
timestamp 1644511149
transform 1 0 57040 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_1_620
timestamp 1644511149
transform 1 0 58144 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_624
timestamp 1644511149
transform 1 0 58512 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_3
timestamp 1644511149
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_15
timestamp 1644511149
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_27
timestamp 1644511149
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_2_29
timestamp 1644511149
transform 1 0 3772 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_53
timestamp 1644511149
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_2_65
timestamp 1644511149
transform 1 0 7084 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_2_80
timestamp 1644511149
transform 1 0 8464 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_2_85
timestamp 1644511149
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_97
timestamp 1644511149
transform 1 0 10028 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_109
timestamp 1644511149
transform 1 0 11132 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_121
timestamp 1644511149
transform 1 0 12236 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_133
timestamp 1644511149
transform 1 0 13340 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_139
timestamp 1644511149
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_141
timestamp 1644511149
transform 1 0 14076 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_166
timestamp 1644511149
transform 1 0 16376 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_170
timestamp 1644511149
transform 1 0 16744 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_192
timestamp 1644511149
transform 1 0 18768 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_2_197
timestamp 1644511149
transform 1 0 19228 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_2_209
timestamp 1644511149
transform 1 0 20332 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_233
timestamp 1644511149
transform 1 0 22540 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_245
timestamp 1644511149
transform 1 0 23644 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_251
timestamp 1644511149
transform 1 0 24196 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_253
timestamp 1644511149
transform 1 0 24380 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_265
timestamp 1644511149
transform 1 0 25484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_277
timestamp 1644511149
transform 1 0 26588 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_289
timestamp 1644511149
transform 1 0 27692 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_301
timestamp 1644511149
transform 1 0 28796 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_307
timestamp 1644511149
transform 1 0 29348 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_309
timestamp 1644511149
transform 1 0 29532 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_321
timestamp 1644511149
transform 1 0 30636 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_333
timestamp 1644511149
transform 1 0 31740 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_345
timestamp 1644511149
transform 1 0 32844 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_357
timestamp 1644511149
transform 1 0 33948 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_363
timestamp 1644511149
transform 1 0 34500 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_365
timestamp 1644511149
transform 1 0 34684 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_377
timestamp 1644511149
transform 1 0 35788 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_389
timestamp 1644511149
transform 1 0 36892 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_401
timestamp 1644511149
transform 1 0 37996 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_413
timestamp 1644511149
transform 1 0 39100 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_419
timestamp 1644511149
transform 1 0 39652 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_421
timestamp 1644511149
transform 1 0 39836 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_433
timestamp 1644511149
transform 1 0 40940 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_445
timestamp 1644511149
transform 1 0 42044 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_457
timestamp 1644511149
transform 1 0 43148 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_472
timestamp 1644511149
transform 1 0 44528 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_2_498
timestamp 1644511149
transform 1 0 46920 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_510
timestamp 1644511149
transform 1 0 48024 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_522
timestamp 1644511149
transform 1 0 49128 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_530
timestamp 1644511149
transform 1 0 49864 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_2_533
timestamp 1644511149
transform 1 0 50140 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_2_545
timestamp 1644511149
transform 1 0 51244 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_569
timestamp 1644511149
transform 1 0 53452 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_584
timestamp 1644511149
transform 1 0 54832 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_589
timestamp 1644511149
transform 1 0 55292 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_596
timestamp 1644511149
transform 1 0 55936 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_621
timestamp 1644511149
transform 1 0 58236 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_3
timestamp 1644511149
transform 1 0 1380 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_3_30
timestamp 1644511149
transform 1 0 3864 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_3_37
timestamp 1644511149
transform 1 0 4508 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_49
timestamp 1644511149
transform 1 0 5612 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_55
timestamp 1644511149
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_57
timestamp 1644511149
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_3_69
timestamp 1644511149
transform 1 0 7452 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_86
timestamp 1644511149
transform 1 0 9016 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_98
timestamp 1644511149
transform 1 0 10120 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_3_110
timestamp 1644511149
transform 1 0 11224 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_3_113
timestamp 1644511149
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_125
timestamp 1644511149
transform 1 0 12604 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_137
timestamp 1644511149
transform 1 0 13708 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_149
timestamp 1644511149
transform 1 0 14812 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_161
timestamp 1644511149
transform 1 0 15916 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_167
timestamp 1644511149
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_169
timestamp 1644511149
transform 1 0 16652 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_181
timestamp 1644511149
transform 1 0 17756 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_193
timestamp 1644511149
transform 1 0 18860 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_205
timestamp 1644511149
transform 1 0 19964 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_3_216
timestamp 1644511149
transform 1 0 20976 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_3_225
timestamp 1644511149
transform 1 0 21804 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_237
timestamp 1644511149
transform 1 0 22908 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_249
timestamp 1644511149
transform 1 0 24012 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_261
timestamp 1644511149
transform 1 0 25116 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_273
timestamp 1644511149
transform 1 0 26220 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_279
timestamp 1644511149
transform 1 0 26772 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_281
timestamp 1644511149
transform 1 0 26956 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_293
timestamp 1644511149
transform 1 0 28060 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_305
timestamp 1644511149
transform 1 0 29164 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_317
timestamp 1644511149
transform 1 0 30268 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_329
timestamp 1644511149
transform 1 0 31372 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_335
timestamp 1644511149
transform 1 0 31924 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_337
timestamp 1644511149
transform 1 0 32108 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_349
timestamp 1644511149
transform 1 0 33212 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_361
timestamp 1644511149
transform 1 0 34316 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_373
timestamp 1644511149
transform 1 0 35420 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_385
timestamp 1644511149
transform 1 0 36524 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_391
timestamp 1644511149
transform 1 0 37076 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_393
timestamp 1644511149
transform 1 0 37260 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_405
timestamp 1644511149
transform 1 0 38364 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_417
timestamp 1644511149
transform 1 0 39468 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_429
timestamp 1644511149
transform 1 0 40572 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_441
timestamp 1644511149
transform 1 0 41676 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_447
timestamp 1644511149
transform 1 0 42228 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_449
timestamp 1644511149
transform 1 0 42412 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_461
timestamp 1644511149
transform 1 0 43516 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_473
timestamp 1644511149
transform 1 0 44620 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_485
timestamp 1644511149
transform 1 0 45724 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_497
timestamp 1644511149
transform 1 0 46828 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_503
timestamp 1644511149
transform 1 0 47380 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_505
timestamp 1644511149
transform 1 0 47564 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_517
timestamp 1644511149
transform 1 0 48668 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_529
timestamp 1644511149
transform 1 0 49772 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_541
timestamp 1644511149
transform 1 0 50876 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_547
timestamp 1644511149
transform 1 0 51428 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_551
timestamp 1644511149
transform 1 0 51796 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_559
timestamp 1644511149
transform 1 0 52532 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_561
timestamp 1644511149
transform 1 0 52716 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_573
timestamp 1644511149
transform 1 0 53820 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_579
timestamp 1644511149
transform 1 0 54372 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_583
timestamp 1644511149
transform 1 0 54740 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_3_612
timestamp 1644511149
transform 1 0 57408 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_620
timestamp 1644511149
transform 1 0 58144 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_624
timestamp 1644511149
transform 1 0 58512 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_3
timestamp 1644511149
transform 1 0 1380 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_11
timestamp 1644511149
transform 1 0 2116 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_4_16
timestamp 1644511149
transform 1 0 2576 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_29
timestamp 1644511149
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_41
timestamp 1644511149
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_53
timestamp 1644511149
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_65
timestamp 1644511149
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_77
timestamp 1644511149
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_83
timestamp 1644511149
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_85
timestamp 1644511149
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_97
timestamp 1644511149
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_109
timestamp 1644511149
transform 1 0 11132 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_121
timestamp 1644511149
transform 1 0 12236 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_133
timestamp 1644511149
transform 1 0 13340 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_139
timestamp 1644511149
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_141
timestamp 1644511149
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_153
timestamp 1644511149
transform 1 0 15180 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_165
timestamp 1644511149
transform 1 0 16284 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_177
timestamp 1644511149
transform 1 0 17388 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_189
timestamp 1644511149
transform 1 0 18492 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_195
timestamp 1644511149
transform 1 0 19044 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_197
timestamp 1644511149
transform 1 0 19228 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_209
timestamp 1644511149
transform 1 0 20332 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_221
timestamp 1644511149
transform 1 0 21436 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_233
timestamp 1644511149
transform 1 0 22540 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_245
timestamp 1644511149
transform 1 0 23644 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_251
timestamp 1644511149
transform 1 0 24196 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_253
timestamp 1644511149
transform 1 0 24380 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_265
timestamp 1644511149
transform 1 0 25484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_277
timestamp 1644511149
transform 1 0 26588 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_289
timestamp 1644511149
transform 1 0 27692 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_301
timestamp 1644511149
transform 1 0 28796 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_307
timestamp 1644511149
transform 1 0 29348 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_309
timestamp 1644511149
transform 1 0 29532 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_321
timestamp 1644511149
transform 1 0 30636 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_333
timestamp 1644511149
transform 1 0 31740 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_345
timestamp 1644511149
transform 1 0 32844 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_357
timestamp 1644511149
transform 1 0 33948 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_363
timestamp 1644511149
transform 1 0 34500 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_365
timestamp 1644511149
transform 1 0 34684 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_377
timestamp 1644511149
transform 1 0 35788 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_389
timestamp 1644511149
transform 1 0 36892 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_401
timestamp 1644511149
transform 1 0 37996 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_413
timestamp 1644511149
transform 1 0 39100 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_419
timestamp 1644511149
transform 1 0 39652 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_421
timestamp 1644511149
transform 1 0 39836 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_433
timestamp 1644511149
transform 1 0 40940 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_445
timestamp 1644511149
transform 1 0 42044 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_457
timestamp 1644511149
transform 1 0 43148 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_469
timestamp 1644511149
transform 1 0 44252 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_475
timestamp 1644511149
transform 1 0 44804 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_477
timestamp 1644511149
transform 1 0 44988 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_489
timestamp 1644511149
transform 1 0 46092 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_501
timestamp 1644511149
transform 1 0 47196 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_513
timestamp 1644511149
transform 1 0 48300 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_525
timestamp 1644511149
transform 1 0 49404 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_531
timestamp 1644511149
transform 1 0 49956 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_533
timestamp 1644511149
transform 1 0 50140 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_545
timestamp 1644511149
transform 1 0 51244 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_557
timestamp 1644511149
transform 1 0 52348 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_569
timestamp 1644511149
transform 1 0 53452 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_581
timestamp 1644511149
transform 1 0 54556 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_587
timestamp 1644511149
transform 1 0 55108 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_589
timestamp 1644511149
transform 1 0 55292 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_4_597
timestamp 1644511149
transform 1 0 56028 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_4_621
timestamp 1644511149
transform 1 0 58236 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_5_3
timestamp 1644511149
transform 1 0 1380 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_9
timestamp 1644511149
transform 1 0 1932 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_13
timestamp 1644511149
transform 1 0 2300 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_25
timestamp 1644511149
transform 1 0 3404 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_37
timestamp 1644511149
transform 1 0 4508 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_49
timestamp 1644511149
transform 1 0 5612 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_55
timestamp 1644511149
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_57
timestamp 1644511149
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_69
timestamp 1644511149
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_81
timestamp 1644511149
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_93
timestamp 1644511149
transform 1 0 9660 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_105
timestamp 1644511149
transform 1 0 10764 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_111
timestamp 1644511149
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_113
timestamp 1644511149
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_125
timestamp 1644511149
transform 1 0 12604 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_137
timestamp 1644511149
transform 1 0 13708 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_149
timestamp 1644511149
transform 1 0 14812 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_161
timestamp 1644511149
transform 1 0 15916 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_167
timestamp 1644511149
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_169
timestamp 1644511149
transform 1 0 16652 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_181
timestamp 1644511149
transform 1 0 17756 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_193
timestamp 1644511149
transform 1 0 18860 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_205
timestamp 1644511149
transform 1 0 19964 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_217
timestamp 1644511149
transform 1 0 21068 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_223
timestamp 1644511149
transform 1 0 21620 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_225
timestamp 1644511149
transform 1 0 21804 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_237
timestamp 1644511149
transform 1 0 22908 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_249
timestamp 1644511149
transform 1 0 24012 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_261
timestamp 1644511149
transform 1 0 25116 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_273
timestamp 1644511149
transform 1 0 26220 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_279
timestamp 1644511149
transform 1 0 26772 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_281
timestamp 1644511149
transform 1 0 26956 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_293
timestamp 1644511149
transform 1 0 28060 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_305
timestamp 1644511149
transform 1 0 29164 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_317
timestamp 1644511149
transform 1 0 30268 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_329
timestamp 1644511149
transform 1 0 31372 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_335
timestamp 1644511149
transform 1 0 31924 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_337
timestamp 1644511149
transform 1 0 32108 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_349
timestamp 1644511149
transform 1 0 33212 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_361
timestamp 1644511149
transform 1 0 34316 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_373
timestamp 1644511149
transform 1 0 35420 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_385
timestamp 1644511149
transform 1 0 36524 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_391
timestamp 1644511149
transform 1 0 37076 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_393
timestamp 1644511149
transform 1 0 37260 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_405
timestamp 1644511149
transform 1 0 38364 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_417
timestamp 1644511149
transform 1 0 39468 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_429
timestamp 1644511149
transform 1 0 40572 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_441
timestamp 1644511149
transform 1 0 41676 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_447
timestamp 1644511149
transform 1 0 42228 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_449
timestamp 1644511149
transform 1 0 42412 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_461
timestamp 1644511149
transform 1 0 43516 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_473
timestamp 1644511149
transform 1 0 44620 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_485
timestamp 1644511149
transform 1 0 45724 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_497
timestamp 1644511149
transform 1 0 46828 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_503
timestamp 1644511149
transform 1 0 47380 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_505
timestamp 1644511149
transform 1 0 47564 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_517
timestamp 1644511149
transform 1 0 48668 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_529
timestamp 1644511149
transform 1 0 49772 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_541
timestamp 1644511149
transform 1 0 50876 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_553
timestamp 1644511149
transform 1 0 51980 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_559
timestamp 1644511149
transform 1 0 52532 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_561
timestamp 1644511149
transform 1 0 52716 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_573
timestamp 1644511149
transform 1 0 53820 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_585
timestamp 1644511149
transform 1 0 54924 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_597
timestamp 1644511149
transform 1 0 56028 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_609
timestamp 1644511149
transform 1 0 57132 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_615
timestamp 1644511149
transform 1 0 57684 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_617
timestamp 1644511149
transform 1 0 57868 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_6_3
timestamp 1644511149
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_15
timestamp 1644511149
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 1644511149
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_29
timestamp 1644511149
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_41
timestamp 1644511149
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_53
timestamp 1644511149
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_65
timestamp 1644511149
transform 1 0 7084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_77
timestamp 1644511149
transform 1 0 8188 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_83
timestamp 1644511149
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_85
timestamp 1644511149
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_97
timestamp 1644511149
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_109
timestamp 1644511149
transform 1 0 11132 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_121
timestamp 1644511149
transform 1 0 12236 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_133
timestamp 1644511149
transform 1 0 13340 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_139
timestamp 1644511149
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_141
timestamp 1644511149
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_153
timestamp 1644511149
transform 1 0 15180 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_165
timestamp 1644511149
transform 1 0 16284 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_177
timestamp 1644511149
transform 1 0 17388 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_189
timestamp 1644511149
transform 1 0 18492 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_195
timestamp 1644511149
transform 1 0 19044 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_197
timestamp 1644511149
transform 1 0 19228 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_209
timestamp 1644511149
transform 1 0 20332 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_221
timestamp 1644511149
transform 1 0 21436 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_233
timestamp 1644511149
transform 1 0 22540 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_245
timestamp 1644511149
transform 1 0 23644 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_251
timestamp 1644511149
transform 1 0 24196 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_253
timestamp 1644511149
transform 1 0 24380 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_265
timestamp 1644511149
transform 1 0 25484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_277
timestamp 1644511149
transform 1 0 26588 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_289
timestamp 1644511149
transform 1 0 27692 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_301
timestamp 1644511149
transform 1 0 28796 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_307
timestamp 1644511149
transform 1 0 29348 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_309
timestamp 1644511149
transform 1 0 29532 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_321
timestamp 1644511149
transform 1 0 30636 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_333
timestamp 1644511149
transform 1 0 31740 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_345
timestamp 1644511149
transform 1 0 32844 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_357
timestamp 1644511149
transform 1 0 33948 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_363
timestamp 1644511149
transform 1 0 34500 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_365
timestamp 1644511149
transform 1 0 34684 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_377
timestamp 1644511149
transform 1 0 35788 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_389
timestamp 1644511149
transform 1 0 36892 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_401
timestamp 1644511149
transform 1 0 37996 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_413
timestamp 1644511149
transform 1 0 39100 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_419
timestamp 1644511149
transform 1 0 39652 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_421
timestamp 1644511149
transform 1 0 39836 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_433
timestamp 1644511149
transform 1 0 40940 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_445
timestamp 1644511149
transform 1 0 42044 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_457
timestamp 1644511149
transform 1 0 43148 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_469
timestamp 1644511149
transform 1 0 44252 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_475
timestamp 1644511149
transform 1 0 44804 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_477
timestamp 1644511149
transform 1 0 44988 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_489
timestamp 1644511149
transform 1 0 46092 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_501
timestamp 1644511149
transform 1 0 47196 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_513
timestamp 1644511149
transform 1 0 48300 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_525
timestamp 1644511149
transform 1 0 49404 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_531
timestamp 1644511149
transform 1 0 49956 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_533
timestamp 1644511149
transform 1 0 50140 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_545
timestamp 1644511149
transform 1 0 51244 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_557
timestamp 1644511149
transform 1 0 52348 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_569
timestamp 1644511149
transform 1 0 53452 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_581
timestamp 1644511149
transform 1 0 54556 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_587
timestamp 1644511149
transform 1 0 55108 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_589
timestamp 1644511149
transform 1 0 55292 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_601
timestamp 1644511149
transform 1 0 56396 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_613
timestamp 1644511149
transform 1 0 57500 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_3
timestamp 1644511149
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_15
timestamp 1644511149
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_27
timestamp 1644511149
transform 1 0 3588 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_39
timestamp 1644511149
transform 1 0 4692 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_51
timestamp 1644511149
transform 1 0 5796 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_55
timestamp 1644511149
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_57
timestamp 1644511149
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_69
timestamp 1644511149
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_81
timestamp 1644511149
transform 1 0 8556 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_93
timestamp 1644511149
transform 1 0 9660 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_105
timestamp 1644511149
transform 1 0 10764 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_111
timestamp 1644511149
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_113
timestamp 1644511149
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_125
timestamp 1644511149
transform 1 0 12604 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_137
timestamp 1644511149
transform 1 0 13708 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_149
timestamp 1644511149
transform 1 0 14812 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_161
timestamp 1644511149
transform 1 0 15916 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_167
timestamp 1644511149
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_169
timestamp 1644511149
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_181
timestamp 1644511149
transform 1 0 17756 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_193
timestamp 1644511149
transform 1 0 18860 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_205
timestamp 1644511149
transform 1 0 19964 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_217
timestamp 1644511149
transform 1 0 21068 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_223
timestamp 1644511149
transform 1 0 21620 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_225
timestamp 1644511149
transform 1 0 21804 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_237
timestamp 1644511149
transform 1 0 22908 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_249
timestamp 1644511149
transform 1 0 24012 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_261
timestamp 1644511149
transform 1 0 25116 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_273
timestamp 1644511149
transform 1 0 26220 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_279
timestamp 1644511149
transform 1 0 26772 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_281
timestamp 1644511149
transform 1 0 26956 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_293
timestamp 1644511149
transform 1 0 28060 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_305
timestamp 1644511149
transform 1 0 29164 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_317
timestamp 1644511149
transform 1 0 30268 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_329
timestamp 1644511149
transform 1 0 31372 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_335
timestamp 1644511149
transform 1 0 31924 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_337
timestamp 1644511149
transform 1 0 32108 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_349
timestamp 1644511149
transform 1 0 33212 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_361
timestamp 1644511149
transform 1 0 34316 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_373
timestamp 1644511149
transform 1 0 35420 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_385
timestamp 1644511149
transform 1 0 36524 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_391
timestamp 1644511149
transform 1 0 37076 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_393
timestamp 1644511149
transform 1 0 37260 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_405
timestamp 1644511149
transform 1 0 38364 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_417
timestamp 1644511149
transform 1 0 39468 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_429
timestamp 1644511149
transform 1 0 40572 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_441
timestamp 1644511149
transform 1 0 41676 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_447
timestamp 1644511149
transform 1 0 42228 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_449
timestamp 1644511149
transform 1 0 42412 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_461
timestamp 1644511149
transform 1 0 43516 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_473
timestamp 1644511149
transform 1 0 44620 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_485
timestamp 1644511149
transform 1 0 45724 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_497
timestamp 1644511149
transform 1 0 46828 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_503
timestamp 1644511149
transform 1 0 47380 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_505
timestamp 1644511149
transform 1 0 47564 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_517
timestamp 1644511149
transform 1 0 48668 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_529
timestamp 1644511149
transform 1 0 49772 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_541
timestamp 1644511149
transform 1 0 50876 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_553
timestamp 1644511149
transform 1 0 51980 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_559
timestamp 1644511149
transform 1 0 52532 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_561
timestamp 1644511149
transform 1 0 52716 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_573
timestamp 1644511149
transform 1 0 53820 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_585
timestamp 1644511149
transform 1 0 54924 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_597
timestamp 1644511149
transform 1 0 56028 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_609
timestamp 1644511149
transform 1 0 57132 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_615
timestamp 1644511149
transform 1 0 57684 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_617
timestamp 1644511149
transform 1 0 57868 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_8_3
timestamp 1644511149
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_15
timestamp 1644511149
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 1644511149
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_29
timestamp 1644511149
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_41
timestamp 1644511149
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_53
timestamp 1644511149
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_65
timestamp 1644511149
transform 1 0 7084 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_77
timestamp 1644511149
transform 1 0 8188 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_83
timestamp 1644511149
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_85
timestamp 1644511149
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_97
timestamp 1644511149
transform 1 0 10028 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_109
timestamp 1644511149
transform 1 0 11132 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_121
timestamp 1644511149
transform 1 0 12236 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_133
timestamp 1644511149
transform 1 0 13340 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_139
timestamp 1644511149
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_141
timestamp 1644511149
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_153
timestamp 1644511149
transform 1 0 15180 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_165
timestamp 1644511149
transform 1 0 16284 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_177
timestamp 1644511149
transform 1 0 17388 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_189
timestamp 1644511149
transform 1 0 18492 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_195
timestamp 1644511149
transform 1 0 19044 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_197
timestamp 1644511149
transform 1 0 19228 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_209
timestamp 1644511149
transform 1 0 20332 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_221
timestamp 1644511149
transform 1 0 21436 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_233
timestamp 1644511149
transform 1 0 22540 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_245
timestamp 1644511149
transform 1 0 23644 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_251
timestamp 1644511149
transform 1 0 24196 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_253
timestamp 1644511149
transform 1 0 24380 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_265
timestamp 1644511149
transform 1 0 25484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_277
timestamp 1644511149
transform 1 0 26588 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_289
timestamp 1644511149
transform 1 0 27692 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_301
timestamp 1644511149
transform 1 0 28796 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_307
timestamp 1644511149
transform 1 0 29348 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_309
timestamp 1644511149
transform 1 0 29532 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_321
timestamp 1644511149
transform 1 0 30636 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_333
timestamp 1644511149
transform 1 0 31740 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_345
timestamp 1644511149
transform 1 0 32844 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_357
timestamp 1644511149
transform 1 0 33948 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_363
timestamp 1644511149
transform 1 0 34500 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_365
timestamp 1644511149
transform 1 0 34684 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_377
timestamp 1644511149
transform 1 0 35788 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_389
timestamp 1644511149
transform 1 0 36892 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_401
timestamp 1644511149
transform 1 0 37996 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_413
timestamp 1644511149
transform 1 0 39100 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_419
timestamp 1644511149
transform 1 0 39652 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_421
timestamp 1644511149
transform 1 0 39836 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_433
timestamp 1644511149
transform 1 0 40940 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_445
timestamp 1644511149
transform 1 0 42044 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_457
timestamp 1644511149
transform 1 0 43148 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_469
timestamp 1644511149
transform 1 0 44252 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_475
timestamp 1644511149
transform 1 0 44804 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_477
timestamp 1644511149
transform 1 0 44988 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_489
timestamp 1644511149
transform 1 0 46092 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_501
timestamp 1644511149
transform 1 0 47196 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_513
timestamp 1644511149
transform 1 0 48300 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_525
timestamp 1644511149
transform 1 0 49404 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_531
timestamp 1644511149
transform 1 0 49956 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_533
timestamp 1644511149
transform 1 0 50140 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_545
timestamp 1644511149
transform 1 0 51244 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_557
timestamp 1644511149
transform 1 0 52348 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_569
timestamp 1644511149
transform 1 0 53452 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_581
timestamp 1644511149
transform 1 0 54556 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_587
timestamp 1644511149
transform 1 0 55108 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_589
timestamp 1644511149
transform 1 0 55292 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_601
timestamp 1644511149
transform 1 0 56396 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_613
timestamp 1644511149
transform 1 0 57500 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_3
timestamp 1644511149
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_15
timestamp 1644511149
transform 1 0 2484 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_27
timestamp 1644511149
transform 1 0 3588 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_39
timestamp 1644511149
transform 1 0 4692 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_51
timestamp 1644511149
transform 1 0 5796 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_55
timestamp 1644511149
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_57
timestamp 1644511149
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_69
timestamp 1644511149
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_81
timestamp 1644511149
transform 1 0 8556 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_93
timestamp 1644511149
transform 1 0 9660 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_105
timestamp 1644511149
transform 1 0 10764 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_111
timestamp 1644511149
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_113
timestamp 1644511149
transform 1 0 11500 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_125
timestamp 1644511149
transform 1 0 12604 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_137
timestamp 1644511149
transform 1 0 13708 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_149
timestamp 1644511149
transform 1 0 14812 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_161
timestamp 1644511149
transform 1 0 15916 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_167
timestamp 1644511149
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_169
timestamp 1644511149
transform 1 0 16652 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_181
timestamp 1644511149
transform 1 0 17756 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_193
timestamp 1644511149
transform 1 0 18860 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_205
timestamp 1644511149
transform 1 0 19964 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_217
timestamp 1644511149
transform 1 0 21068 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_223
timestamp 1644511149
transform 1 0 21620 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_225
timestamp 1644511149
transform 1 0 21804 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_237
timestamp 1644511149
transform 1 0 22908 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_249
timestamp 1644511149
transform 1 0 24012 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_261
timestamp 1644511149
transform 1 0 25116 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_273
timestamp 1644511149
transform 1 0 26220 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_279
timestamp 1644511149
transform 1 0 26772 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_281
timestamp 1644511149
transform 1 0 26956 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_293
timestamp 1644511149
transform 1 0 28060 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_305
timestamp 1644511149
transform 1 0 29164 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_317
timestamp 1644511149
transform 1 0 30268 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_329
timestamp 1644511149
transform 1 0 31372 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_335
timestamp 1644511149
transform 1 0 31924 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_337
timestamp 1644511149
transform 1 0 32108 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_349
timestamp 1644511149
transform 1 0 33212 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_361
timestamp 1644511149
transform 1 0 34316 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_373
timestamp 1644511149
transform 1 0 35420 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_385
timestamp 1644511149
transform 1 0 36524 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_391
timestamp 1644511149
transform 1 0 37076 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_393
timestamp 1644511149
transform 1 0 37260 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_405
timestamp 1644511149
transform 1 0 38364 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_417
timestamp 1644511149
transform 1 0 39468 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_429
timestamp 1644511149
transform 1 0 40572 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_441
timestamp 1644511149
transform 1 0 41676 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_447
timestamp 1644511149
transform 1 0 42228 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_449
timestamp 1644511149
transform 1 0 42412 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_461
timestamp 1644511149
transform 1 0 43516 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_473
timestamp 1644511149
transform 1 0 44620 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_485
timestamp 1644511149
transform 1 0 45724 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_497
timestamp 1644511149
transform 1 0 46828 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_503
timestamp 1644511149
transform 1 0 47380 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_505
timestamp 1644511149
transform 1 0 47564 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_517
timestamp 1644511149
transform 1 0 48668 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_529
timestamp 1644511149
transform 1 0 49772 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_541
timestamp 1644511149
transform 1 0 50876 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_553
timestamp 1644511149
transform 1 0 51980 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_559
timestamp 1644511149
transform 1 0 52532 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_561
timestamp 1644511149
transform 1 0 52716 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_573
timestamp 1644511149
transform 1 0 53820 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_585
timestamp 1644511149
transform 1 0 54924 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_597
timestamp 1644511149
transform 1 0 56028 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_609
timestamp 1644511149
transform 1 0 57132 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_615
timestamp 1644511149
transform 1 0 57684 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_617
timestamp 1644511149
transform 1 0 57868 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_10_3
timestamp 1644511149
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_15
timestamp 1644511149
transform 1 0 2484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp 1644511149
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_29
timestamp 1644511149
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_41
timestamp 1644511149
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_53
timestamp 1644511149
transform 1 0 5980 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_65
timestamp 1644511149
transform 1 0 7084 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_77
timestamp 1644511149
transform 1 0 8188 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_83
timestamp 1644511149
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_85
timestamp 1644511149
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_97
timestamp 1644511149
transform 1 0 10028 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_109
timestamp 1644511149
transform 1 0 11132 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_121
timestamp 1644511149
transform 1 0 12236 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_133
timestamp 1644511149
transform 1 0 13340 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_139
timestamp 1644511149
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_141
timestamp 1644511149
transform 1 0 14076 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_153
timestamp 1644511149
transform 1 0 15180 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_165
timestamp 1644511149
transform 1 0 16284 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_177
timestamp 1644511149
transform 1 0 17388 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_189
timestamp 1644511149
transform 1 0 18492 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_195
timestamp 1644511149
transform 1 0 19044 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_197
timestamp 1644511149
transform 1 0 19228 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_209
timestamp 1644511149
transform 1 0 20332 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_221
timestamp 1644511149
transform 1 0 21436 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_233
timestamp 1644511149
transform 1 0 22540 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_245
timestamp 1644511149
transform 1 0 23644 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_251
timestamp 1644511149
transform 1 0 24196 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_253
timestamp 1644511149
transform 1 0 24380 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_265
timestamp 1644511149
transform 1 0 25484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_277
timestamp 1644511149
transform 1 0 26588 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_289
timestamp 1644511149
transform 1 0 27692 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_301
timestamp 1644511149
transform 1 0 28796 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_307
timestamp 1644511149
transform 1 0 29348 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_309
timestamp 1644511149
transform 1 0 29532 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_321
timestamp 1644511149
transform 1 0 30636 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_333
timestamp 1644511149
transform 1 0 31740 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_345
timestamp 1644511149
transform 1 0 32844 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_357
timestamp 1644511149
transform 1 0 33948 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_363
timestamp 1644511149
transform 1 0 34500 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_365
timestamp 1644511149
transform 1 0 34684 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_377
timestamp 1644511149
transform 1 0 35788 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_389
timestamp 1644511149
transform 1 0 36892 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_401
timestamp 1644511149
transform 1 0 37996 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_413
timestamp 1644511149
transform 1 0 39100 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_419
timestamp 1644511149
transform 1 0 39652 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_421
timestamp 1644511149
transform 1 0 39836 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_433
timestamp 1644511149
transform 1 0 40940 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_445
timestamp 1644511149
transform 1 0 42044 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_457
timestamp 1644511149
transform 1 0 43148 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_469
timestamp 1644511149
transform 1 0 44252 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_475
timestamp 1644511149
transform 1 0 44804 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_477
timestamp 1644511149
transform 1 0 44988 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_489
timestamp 1644511149
transform 1 0 46092 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_501
timestamp 1644511149
transform 1 0 47196 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_513
timestamp 1644511149
transform 1 0 48300 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_525
timestamp 1644511149
transform 1 0 49404 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_531
timestamp 1644511149
transform 1 0 49956 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_533
timestamp 1644511149
transform 1 0 50140 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_545
timestamp 1644511149
transform 1 0 51244 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_557
timestamp 1644511149
transform 1 0 52348 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_569
timestamp 1644511149
transform 1 0 53452 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_581
timestamp 1644511149
transform 1 0 54556 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_587
timestamp 1644511149
transform 1 0 55108 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_589
timestamp 1644511149
transform 1 0 55292 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_601
timestamp 1644511149
transform 1 0 56396 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_613
timestamp 1644511149
transform 1 0 57500 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_3
timestamp 1644511149
transform 1 0 1380 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_15
timestamp 1644511149
transform 1 0 2484 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_27
timestamp 1644511149
transform 1 0 3588 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_39
timestamp 1644511149
transform 1 0 4692 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_51
timestamp 1644511149
transform 1 0 5796 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_55
timestamp 1644511149
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_57
timestamp 1644511149
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_69
timestamp 1644511149
transform 1 0 7452 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_81
timestamp 1644511149
transform 1 0 8556 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_93
timestamp 1644511149
transform 1 0 9660 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_105
timestamp 1644511149
transform 1 0 10764 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_111
timestamp 1644511149
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_113
timestamp 1644511149
transform 1 0 11500 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_125
timestamp 1644511149
transform 1 0 12604 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_137
timestamp 1644511149
transform 1 0 13708 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_149
timestamp 1644511149
transform 1 0 14812 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_161
timestamp 1644511149
transform 1 0 15916 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_167
timestamp 1644511149
transform 1 0 16468 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_169
timestamp 1644511149
transform 1 0 16652 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_181
timestamp 1644511149
transform 1 0 17756 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_193
timestamp 1644511149
transform 1 0 18860 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_205
timestamp 1644511149
transform 1 0 19964 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_217
timestamp 1644511149
transform 1 0 21068 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_223
timestamp 1644511149
transform 1 0 21620 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_225
timestamp 1644511149
transform 1 0 21804 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_237
timestamp 1644511149
transform 1 0 22908 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_249
timestamp 1644511149
transform 1 0 24012 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_261
timestamp 1644511149
transform 1 0 25116 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_273
timestamp 1644511149
transform 1 0 26220 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_279
timestamp 1644511149
transform 1 0 26772 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_281
timestamp 1644511149
transform 1 0 26956 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_293
timestamp 1644511149
transform 1 0 28060 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_305
timestamp 1644511149
transform 1 0 29164 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_317
timestamp 1644511149
transform 1 0 30268 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_329
timestamp 1644511149
transform 1 0 31372 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_335
timestamp 1644511149
transform 1 0 31924 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_337
timestamp 1644511149
transform 1 0 32108 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_349
timestamp 1644511149
transform 1 0 33212 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_361
timestamp 1644511149
transform 1 0 34316 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_373
timestamp 1644511149
transform 1 0 35420 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_385
timestamp 1644511149
transform 1 0 36524 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_391
timestamp 1644511149
transform 1 0 37076 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_393
timestamp 1644511149
transform 1 0 37260 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_405
timestamp 1644511149
transform 1 0 38364 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_417
timestamp 1644511149
transform 1 0 39468 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_429
timestamp 1644511149
transform 1 0 40572 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_441
timestamp 1644511149
transform 1 0 41676 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_447
timestamp 1644511149
transform 1 0 42228 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_449
timestamp 1644511149
transform 1 0 42412 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_461
timestamp 1644511149
transform 1 0 43516 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_473
timestamp 1644511149
transform 1 0 44620 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_485
timestamp 1644511149
transform 1 0 45724 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_497
timestamp 1644511149
transform 1 0 46828 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_503
timestamp 1644511149
transform 1 0 47380 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_505
timestamp 1644511149
transform 1 0 47564 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_517
timestamp 1644511149
transform 1 0 48668 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_529
timestamp 1644511149
transform 1 0 49772 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_541
timestamp 1644511149
transform 1 0 50876 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_553
timestamp 1644511149
transform 1 0 51980 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_559
timestamp 1644511149
transform 1 0 52532 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_561
timestamp 1644511149
transform 1 0 52716 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_573
timestamp 1644511149
transform 1 0 53820 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_585
timestamp 1644511149
transform 1 0 54924 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_11_597
timestamp 1644511149
transform 1 0 56028 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_11_603
timestamp 1644511149
transform 1 0 56580 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_11_615
timestamp 1644511149
transform 1 0 57684 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_620
timestamp 1644511149
transform 1 0 58144 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_624
timestamp 1644511149
transform 1 0 58512 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_3
timestamp 1644511149
transform 1 0 1380 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_15
timestamp 1644511149
transform 1 0 2484 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_27
timestamp 1644511149
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_29
timestamp 1644511149
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_41
timestamp 1644511149
transform 1 0 4876 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_53
timestamp 1644511149
transform 1 0 5980 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_65
timestamp 1644511149
transform 1 0 7084 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_77
timestamp 1644511149
transform 1 0 8188 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_83
timestamp 1644511149
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_85
timestamp 1644511149
transform 1 0 8924 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_97
timestamp 1644511149
transform 1 0 10028 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_109
timestamp 1644511149
transform 1 0 11132 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_121
timestamp 1644511149
transform 1 0 12236 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_133
timestamp 1644511149
transform 1 0 13340 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_139
timestamp 1644511149
transform 1 0 13892 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_141
timestamp 1644511149
transform 1 0 14076 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_153
timestamp 1644511149
transform 1 0 15180 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_165
timestamp 1644511149
transform 1 0 16284 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_177
timestamp 1644511149
transform 1 0 17388 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_189
timestamp 1644511149
transform 1 0 18492 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_195
timestamp 1644511149
transform 1 0 19044 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_197
timestamp 1644511149
transform 1 0 19228 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_209
timestamp 1644511149
transform 1 0 20332 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_221
timestamp 1644511149
transform 1 0 21436 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_233
timestamp 1644511149
transform 1 0 22540 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_245
timestamp 1644511149
transform 1 0 23644 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_251
timestamp 1644511149
transform 1 0 24196 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_253
timestamp 1644511149
transform 1 0 24380 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_265
timestamp 1644511149
transform 1 0 25484 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_277
timestamp 1644511149
transform 1 0 26588 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_289
timestamp 1644511149
transform 1 0 27692 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_301
timestamp 1644511149
transform 1 0 28796 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_307
timestamp 1644511149
transform 1 0 29348 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_309
timestamp 1644511149
transform 1 0 29532 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_321
timestamp 1644511149
transform 1 0 30636 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_333
timestamp 1644511149
transform 1 0 31740 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_345
timestamp 1644511149
transform 1 0 32844 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_357
timestamp 1644511149
transform 1 0 33948 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_363
timestamp 1644511149
transform 1 0 34500 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_365
timestamp 1644511149
transform 1 0 34684 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_377
timestamp 1644511149
transform 1 0 35788 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_389
timestamp 1644511149
transform 1 0 36892 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_401
timestamp 1644511149
transform 1 0 37996 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_413
timestamp 1644511149
transform 1 0 39100 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_419
timestamp 1644511149
transform 1 0 39652 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_421
timestamp 1644511149
transform 1 0 39836 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_433
timestamp 1644511149
transform 1 0 40940 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_445
timestamp 1644511149
transform 1 0 42044 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_457
timestamp 1644511149
transform 1 0 43148 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_469
timestamp 1644511149
transform 1 0 44252 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_475
timestamp 1644511149
transform 1 0 44804 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_477
timestamp 1644511149
transform 1 0 44988 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_489
timestamp 1644511149
transform 1 0 46092 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_501
timestamp 1644511149
transform 1 0 47196 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_513
timestamp 1644511149
transform 1 0 48300 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_525
timestamp 1644511149
transform 1 0 49404 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_531
timestamp 1644511149
transform 1 0 49956 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_533
timestamp 1644511149
transform 1 0 50140 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_545
timestamp 1644511149
transform 1 0 51244 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_557
timestamp 1644511149
transform 1 0 52348 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_569
timestamp 1644511149
transform 1 0 53452 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_581
timestamp 1644511149
transform 1 0 54556 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_587
timestamp 1644511149
transform 1 0 55108 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_589
timestamp 1644511149
transform 1 0 55292 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_12_597
timestamp 1644511149
transform 1 0 56028 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_12_621
timestamp 1644511149
transform 1 0 58236 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_13_3
timestamp 1644511149
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_15
timestamp 1644511149
transform 1 0 2484 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_27
timestamp 1644511149
transform 1 0 3588 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_39
timestamp 1644511149
transform 1 0 4692 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_51
timestamp 1644511149
transform 1 0 5796 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_55
timestamp 1644511149
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_57
timestamp 1644511149
transform 1 0 6348 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_69
timestamp 1644511149
transform 1 0 7452 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_81
timestamp 1644511149
transform 1 0 8556 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_93
timestamp 1644511149
transform 1 0 9660 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_105
timestamp 1644511149
transform 1 0 10764 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_111
timestamp 1644511149
transform 1 0 11316 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_113
timestamp 1644511149
transform 1 0 11500 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_125
timestamp 1644511149
transform 1 0 12604 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_137
timestamp 1644511149
transform 1 0 13708 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_149
timestamp 1644511149
transform 1 0 14812 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_161
timestamp 1644511149
transform 1 0 15916 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_167
timestamp 1644511149
transform 1 0 16468 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_169
timestamp 1644511149
transform 1 0 16652 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_181
timestamp 1644511149
transform 1 0 17756 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_193
timestamp 1644511149
transform 1 0 18860 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_205
timestamp 1644511149
transform 1 0 19964 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_217
timestamp 1644511149
transform 1 0 21068 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_223
timestamp 1644511149
transform 1 0 21620 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_225
timestamp 1644511149
transform 1 0 21804 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_237
timestamp 1644511149
transform 1 0 22908 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_249
timestamp 1644511149
transform 1 0 24012 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_261
timestamp 1644511149
transform 1 0 25116 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_273
timestamp 1644511149
transform 1 0 26220 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_279
timestamp 1644511149
transform 1 0 26772 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_281
timestamp 1644511149
transform 1 0 26956 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_293
timestamp 1644511149
transform 1 0 28060 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_305
timestamp 1644511149
transform 1 0 29164 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_317
timestamp 1644511149
transform 1 0 30268 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_329
timestamp 1644511149
transform 1 0 31372 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_335
timestamp 1644511149
transform 1 0 31924 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_337
timestamp 1644511149
transform 1 0 32108 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_349
timestamp 1644511149
transform 1 0 33212 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_361
timestamp 1644511149
transform 1 0 34316 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_373
timestamp 1644511149
transform 1 0 35420 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_385
timestamp 1644511149
transform 1 0 36524 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_391
timestamp 1644511149
transform 1 0 37076 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_393
timestamp 1644511149
transform 1 0 37260 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_405
timestamp 1644511149
transform 1 0 38364 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_417
timestamp 1644511149
transform 1 0 39468 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_429
timestamp 1644511149
transform 1 0 40572 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_441
timestamp 1644511149
transform 1 0 41676 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_447
timestamp 1644511149
transform 1 0 42228 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_449
timestamp 1644511149
transform 1 0 42412 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_461
timestamp 1644511149
transform 1 0 43516 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_473
timestamp 1644511149
transform 1 0 44620 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_485
timestamp 1644511149
transform 1 0 45724 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_497
timestamp 1644511149
transform 1 0 46828 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_503
timestamp 1644511149
transform 1 0 47380 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_505
timestamp 1644511149
transform 1 0 47564 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_517
timestamp 1644511149
transform 1 0 48668 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_529
timestamp 1644511149
transform 1 0 49772 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_541
timestamp 1644511149
transform 1 0 50876 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_553
timestamp 1644511149
transform 1 0 51980 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_559
timestamp 1644511149
transform 1 0 52532 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_561
timestamp 1644511149
transform 1 0 52716 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_573
timestamp 1644511149
transform 1 0 53820 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_585
timestamp 1644511149
transform 1 0 54924 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_597
timestamp 1644511149
transform 1 0 56028 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_609
timestamp 1644511149
transform 1 0 57132 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_615
timestamp 1644511149
transform 1 0 57684 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_617
timestamp 1644511149
transform 1 0 57868 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_14_3
timestamp 1644511149
transform 1 0 1380 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_9
timestamp 1644511149
transform 1 0 1932 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_13
timestamp 1644511149
transform 1 0 2300 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_14_25
timestamp 1644511149
transform 1 0 3404 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_14_29
timestamp 1644511149
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_41
timestamp 1644511149
transform 1 0 4876 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_53
timestamp 1644511149
transform 1 0 5980 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_65
timestamp 1644511149
transform 1 0 7084 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_77
timestamp 1644511149
transform 1 0 8188 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_83
timestamp 1644511149
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_85
timestamp 1644511149
transform 1 0 8924 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_97
timestamp 1644511149
transform 1 0 10028 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_109
timestamp 1644511149
transform 1 0 11132 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_121
timestamp 1644511149
transform 1 0 12236 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_133
timestamp 1644511149
transform 1 0 13340 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_139
timestamp 1644511149
transform 1 0 13892 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_141
timestamp 1644511149
transform 1 0 14076 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_153
timestamp 1644511149
transform 1 0 15180 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_165
timestamp 1644511149
transform 1 0 16284 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_177
timestamp 1644511149
transform 1 0 17388 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_189
timestamp 1644511149
transform 1 0 18492 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_195
timestamp 1644511149
transform 1 0 19044 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_197
timestamp 1644511149
transform 1 0 19228 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_209
timestamp 1644511149
transform 1 0 20332 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_221
timestamp 1644511149
transform 1 0 21436 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_233
timestamp 1644511149
transform 1 0 22540 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_245
timestamp 1644511149
transform 1 0 23644 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_251
timestamp 1644511149
transform 1 0 24196 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_253
timestamp 1644511149
transform 1 0 24380 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_265
timestamp 1644511149
transform 1 0 25484 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_277
timestamp 1644511149
transform 1 0 26588 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_289
timestamp 1644511149
transform 1 0 27692 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_301
timestamp 1644511149
transform 1 0 28796 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_307
timestamp 1644511149
transform 1 0 29348 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_309
timestamp 1644511149
transform 1 0 29532 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_321
timestamp 1644511149
transform 1 0 30636 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_333
timestamp 1644511149
transform 1 0 31740 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_345
timestamp 1644511149
transform 1 0 32844 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_357
timestamp 1644511149
transform 1 0 33948 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_363
timestamp 1644511149
transform 1 0 34500 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_365
timestamp 1644511149
transform 1 0 34684 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_377
timestamp 1644511149
transform 1 0 35788 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_389
timestamp 1644511149
transform 1 0 36892 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_401
timestamp 1644511149
transform 1 0 37996 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_413
timestamp 1644511149
transform 1 0 39100 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_419
timestamp 1644511149
transform 1 0 39652 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_421
timestamp 1644511149
transform 1 0 39836 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_433
timestamp 1644511149
transform 1 0 40940 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_445
timestamp 1644511149
transform 1 0 42044 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_457
timestamp 1644511149
transform 1 0 43148 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_469
timestamp 1644511149
transform 1 0 44252 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_475
timestamp 1644511149
transform 1 0 44804 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_477
timestamp 1644511149
transform 1 0 44988 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_489
timestamp 1644511149
transform 1 0 46092 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_501
timestamp 1644511149
transform 1 0 47196 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_513
timestamp 1644511149
transform 1 0 48300 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_525
timestamp 1644511149
transform 1 0 49404 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_531
timestamp 1644511149
transform 1 0 49956 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_533
timestamp 1644511149
transform 1 0 50140 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_545
timestamp 1644511149
transform 1 0 51244 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_557
timestamp 1644511149
transform 1 0 52348 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_569
timestamp 1644511149
transform 1 0 53452 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_581
timestamp 1644511149
transform 1 0 54556 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_587
timestamp 1644511149
transform 1 0 55108 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_589
timestamp 1644511149
transform 1 0 55292 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_601
timestamp 1644511149
transform 1 0 56396 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_613
timestamp 1644511149
transform 1 0 57500 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_3
timestamp 1644511149
transform 1 0 1380 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_15_30
timestamp 1644511149
transform 1 0 3864 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_42
timestamp 1644511149
transform 1 0 4968 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_15_54
timestamp 1644511149
transform 1 0 6072 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_15_57
timestamp 1644511149
transform 1 0 6348 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_69
timestamp 1644511149
transform 1 0 7452 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_81
timestamp 1644511149
transform 1 0 8556 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_93
timestamp 1644511149
transform 1 0 9660 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_105
timestamp 1644511149
transform 1 0 10764 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_111
timestamp 1644511149
transform 1 0 11316 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_113
timestamp 1644511149
transform 1 0 11500 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_125
timestamp 1644511149
transform 1 0 12604 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_137
timestamp 1644511149
transform 1 0 13708 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_149
timestamp 1644511149
transform 1 0 14812 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_161
timestamp 1644511149
transform 1 0 15916 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_167
timestamp 1644511149
transform 1 0 16468 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_169
timestamp 1644511149
transform 1 0 16652 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_181
timestamp 1644511149
transform 1 0 17756 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_193
timestamp 1644511149
transform 1 0 18860 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_205
timestamp 1644511149
transform 1 0 19964 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_217
timestamp 1644511149
transform 1 0 21068 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_223
timestamp 1644511149
transform 1 0 21620 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_225
timestamp 1644511149
transform 1 0 21804 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_237
timestamp 1644511149
transform 1 0 22908 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_249
timestamp 1644511149
transform 1 0 24012 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_261
timestamp 1644511149
transform 1 0 25116 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_273
timestamp 1644511149
transform 1 0 26220 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_279
timestamp 1644511149
transform 1 0 26772 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_281
timestamp 1644511149
transform 1 0 26956 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_293
timestamp 1644511149
transform 1 0 28060 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_305
timestamp 1644511149
transform 1 0 29164 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_317
timestamp 1644511149
transform 1 0 30268 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_329
timestamp 1644511149
transform 1 0 31372 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_335
timestamp 1644511149
transform 1 0 31924 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_337
timestamp 1644511149
transform 1 0 32108 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_349
timestamp 1644511149
transform 1 0 33212 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_361
timestamp 1644511149
transform 1 0 34316 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_373
timestamp 1644511149
transform 1 0 35420 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_385
timestamp 1644511149
transform 1 0 36524 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_391
timestamp 1644511149
transform 1 0 37076 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_393
timestamp 1644511149
transform 1 0 37260 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_405
timestamp 1644511149
transform 1 0 38364 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_417
timestamp 1644511149
transform 1 0 39468 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_429
timestamp 1644511149
transform 1 0 40572 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_441
timestamp 1644511149
transform 1 0 41676 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_447
timestamp 1644511149
transform 1 0 42228 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_449
timestamp 1644511149
transform 1 0 42412 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_461
timestamp 1644511149
transform 1 0 43516 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_473
timestamp 1644511149
transform 1 0 44620 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_485
timestamp 1644511149
transform 1 0 45724 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_497
timestamp 1644511149
transform 1 0 46828 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_503
timestamp 1644511149
transform 1 0 47380 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_505
timestamp 1644511149
transform 1 0 47564 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_517
timestamp 1644511149
transform 1 0 48668 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_529
timestamp 1644511149
transform 1 0 49772 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_541
timestamp 1644511149
transform 1 0 50876 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_553
timestamp 1644511149
transform 1 0 51980 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_559
timestamp 1644511149
transform 1 0 52532 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_561
timestamp 1644511149
transform 1 0 52716 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_573
timestamp 1644511149
transform 1 0 53820 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_585
timestamp 1644511149
transform 1 0 54924 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_597
timestamp 1644511149
transform 1 0 56028 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_609
timestamp 1644511149
transform 1 0 57132 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_615
timestamp 1644511149
transform 1 0 57684 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_617
timestamp 1644511149
transform 1 0 57868 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_16_3
timestamp 1644511149
transform 1 0 1380 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_11
timestamp 1644511149
transform 1 0 2116 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_16_16
timestamp 1644511149
transform 1 0 2576 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_29
timestamp 1644511149
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_41
timestamp 1644511149
transform 1 0 4876 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_53
timestamp 1644511149
transform 1 0 5980 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_65
timestamp 1644511149
transform 1 0 7084 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_77
timestamp 1644511149
transform 1 0 8188 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_83
timestamp 1644511149
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_85
timestamp 1644511149
transform 1 0 8924 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_97
timestamp 1644511149
transform 1 0 10028 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_109
timestamp 1644511149
transform 1 0 11132 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_121
timestamp 1644511149
transform 1 0 12236 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_133
timestamp 1644511149
transform 1 0 13340 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_139
timestamp 1644511149
transform 1 0 13892 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_141
timestamp 1644511149
transform 1 0 14076 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_153
timestamp 1644511149
transform 1 0 15180 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_165
timestamp 1644511149
transform 1 0 16284 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_177
timestamp 1644511149
transform 1 0 17388 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_189
timestamp 1644511149
transform 1 0 18492 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_195
timestamp 1644511149
transform 1 0 19044 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_197
timestamp 1644511149
transform 1 0 19228 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_209
timestamp 1644511149
transform 1 0 20332 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_221
timestamp 1644511149
transform 1 0 21436 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_233
timestamp 1644511149
transform 1 0 22540 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_245
timestamp 1644511149
transform 1 0 23644 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_251
timestamp 1644511149
transform 1 0 24196 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_253
timestamp 1644511149
transform 1 0 24380 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_265
timestamp 1644511149
transform 1 0 25484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_277
timestamp 1644511149
transform 1 0 26588 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_289
timestamp 1644511149
transform 1 0 27692 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_301
timestamp 1644511149
transform 1 0 28796 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_307
timestamp 1644511149
transform 1 0 29348 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_309
timestamp 1644511149
transform 1 0 29532 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_321
timestamp 1644511149
transform 1 0 30636 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_333
timestamp 1644511149
transform 1 0 31740 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_345
timestamp 1644511149
transform 1 0 32844 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_357
timestamp 1644511149
transform 1 0 33948 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_363
timestamp 1644511149
transform 1 0 34500 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_365
timestamp 1644511149
transform 1 0 34684 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_377
timestamp 1644511149
transform 1 0 35788 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_389
timestamp 1644511149
transform 1 0 36892 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_401
timestamp 1644511149
transform 1 0 37996 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_413
timestamp 1644511149
transform 1 0 39100 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_419
timestamp 1644511149
transform 1 0 39652 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_421
timestamp 1644511149
transform 1 0 39836 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_433
timestamp 1644511149
transform 1 0 40940 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_445
timestamp 1644511149
transform 1 0 42044 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_457
timestamp 1644511149
transform 1 0 43148 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_469
timestamp 1644511149
transform 1 0 44252 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_475
timestamp 1644511149
transform 1 0 44804 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_477
timestamp 1644511149
transform 1 0 44988 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_489
timestamp 1644511149
transform 1 0 46092 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_501
timestamp 1644511149
transform 1 0 47196 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_513
timestamp 1644511149
transform 1 0 48300 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_525
timestamp 1644511149
transform 1 0 49404 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_531
timestamp 1644511149
transform 1 0 49956 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_533
timestamp 1644511149
transform 1 0 50140 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_545
timestamp 1644511149
transform 1 0 51244 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_557
timestamp 1644511149
transform 1 0 52348 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_569
timestamp 1644511149
transform 1 0 53452 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_581
timestamp 1644511149
transform 1 0 54556 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_587
timestamp 1644511149
transform 1 0 55108 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_589
timestamp 1644511149
transform 1 0 55292 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_16_597
timestamp 1644511149
transform 1 0 56028 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_16_621
timestamp 1644511149
transform 1 0 58236 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_17_3
timestamp 1644511149
transform 1 0 1380 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_15
timestamp 1644511149
transform 1 0 2484 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_27
timestamp 1644511149
transform 1 0 3588 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_39
timestamp 1644511149
transform 1 0 4692 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_51
timestamp 1644511149
transform 1 0 5796 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_55
timestamp 1644511149
transform 1 0 6164 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_57
timestamp 1644511149
transform 1 0 6348 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_69
timestamp 1644511149
transform 1 0 7452 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_81
timestamp 1644511149
transform 1 0 8556 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_93
timestamp 1644511149
transform 1 0 9660 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_105
timestamp 1644511149
transform 1 0 10764 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_111
timestamp 1644511149
transform 1 0 11316 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_113
timestamp 1644511149
transform 1 0 11500 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_125
timestamp 1644511149
transform 1 0 12604 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_137
timestamp 1644511149
transform 1 0 13708 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_149
timestamp 1644511149
transform 1 0 14812 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_161
timestamp 1644511149
transform 1 0 15916 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_167
timestamp 1644511149
transform 1 0 16468 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_169
timestamp 1644511149
transform 1 0 16652 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_181
timestamp 1644511149
transform 1 0 17756 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_193
timestamp 1644511149
transform 1 0 18860 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_205
timestamp 1644511149
transform 1 0 19964 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_217
timestamp 1644511149
transform 1 0 21068 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_223
timestamp 1644511149
transform 1 0 21620 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_225
timestamp 1644511149
transform 1 0 21804 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_237
timestamp 1644511149
transform 1 0 22908 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_249
timestamp 1644511149
transform 1 0 24012 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_261
timestamp 1644511149
transform 1 0 25116 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_273
timestamp 1644511149
transform 1 0 26220 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_279
timestamp 1644511149
transform 1 0 26772 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_281
timestamp 1644511149
transform 1 0 26956 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_293
timestamp 1644511149
transform 1 0 28060 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_305
timestamp 1644511149
transform 1 0 29164 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_317
timestamp 1644511149
transform 1 0 30268 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_329
timestamp 1644511149
transform 1 0 31372 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_335
timestamp 1644511149
transform 1 0 31924 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_337
timestamp 1644511149
transform 1 0 32108 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_349
timestamp 1644511149
transform 1 0 33212 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_361
timestamp 1644511149
transform 1 0 34316 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_373
timestamp 1644511149
transform 1 0 35420 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_385
timestamp 1644511149
transform 1 0 36524 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_391
timestamp 1644511149
transform 1 0 37076 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_393
timestamp 1644511149
transform 1 0 37260 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_405
timestamp 1644511149
transform 1 0 38364 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_417
timestamp 1644511149
transform 1 0 39468 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_429
timestamp 1644511149
transform 1 0 40572 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_441
timestamp 1644511149
transform 1 0 41676 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_447
timestamp 1644511149
transform 1 0 42228 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_449
timestamp 1644511149
transform 1 0 42412 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_461
timestamp 1644511149
transform 1 0 43516 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_473
timestamp 1644511149
transform 1 0 44620 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_485
timestamp 1644511149
transform 1 0 45724 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_497
timestamp 1644511149
transform 1 0 46828 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_503
timestamp 1644511149
transform 1 0 47380 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_505
timestamp 1644511149
transform 1 0 47564 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_517
timestamp 1644511149
transform 1 0 48668 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_529
timestamp 1644511149
transform 1 0 49772 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_541
timestamp 1644511149
transform 1 0 50876 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_553
timestamp 1644511149
transform 1 0 51980 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_559
timestamp 1644511149
transform 1 0 52532 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_561
timestamp 1644511149
transform 1 0 52716 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_573
timestamp 1644511149
transform 1 0 53820 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_585
timestamp 1644511149
transform 1 0 54924 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_597
timestamp 1644511149
transform 1 0 56028 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_605
timestamp 1644511149
transform 1 0 56764 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_17_610
timestamp 1644511149
transform 1 0 57224 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_17_617
timestamp 1644511149
transform 1 0 57868 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_18_3
timestamp 1644511149
transform 1 0 1380 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_15
timestamp 1644511149
transform 1 0 2484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_27
timestamp 1644511149
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_29
timestamp 1644511149
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_41
timestamp 1644511149
transform 1 0 4876 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_53
timestamp 1644511149
transform 1 0 5980 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_65
timestamp 1644511149
transform 1 0 7084 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_77
timestamp 1644511149
transform 1 0 8188 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_83
timestamp 1644511149
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_85
timestamp 1644511149
transform 1 0 8924 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_97
timestamp 1644511149
transform 1 0 10028 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_109
timestamp 1644511149
transform 1 0 11132 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_121
timestamp 1644511149
transform 1 0 12236 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_133
timestamp 1644511149
transform 1 0 13340 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_139
timestamp 1644511149
transform 1 0 13892 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_141
timestamp 1644511149
transform 1 0 14076 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_153
timestamp 1644511149
transform 1 0 15180 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_165
timestamp 1644511149
transform 1 0 16284 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_177
timestamp 1644511149
transform 1 0 17388 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_189
timestamp 1644511149
transform 1 0 18492 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_195
timestamp 1644511149
transform 1 0 19044 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_197
timestamp 1644511149
transform 1 0 19228 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_209
timestamp 1644511149
transform 1 0 20332 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_221
timestamp 1644511149
transform 1 0 21436 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_233
timestamp 1644511149
transform 1 0 22540 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_245
timestamp 1644511149
transform 1 0 23644 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_251
timestamp 1644511149
transform 1 0 24196 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_253
timestamp 1644511149
transform 1 0 24380 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_265
timestamp 1644511149
transform 1 0 25484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_277
timestamp 1644511149
transform 1 0 26588 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_289
timestamp 1644511149
transform 1 0 27692 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_301
timestamp 1644511149
transform 1 0 28796 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_307
timestamp 1644511149
transform 1 0 29348 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_309
timestamp 1644511149
transform 1 0 29532 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_321
timestamp 1644511149
transform 1 0 30636 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_333
timestamp 1644511149
transform 1 0 31740 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_345
timestamp 1644511149
transform 1 0 32844 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_357
timestamp 1644511149
transform 1 0 33948 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_363
timestamp 1644511149
transform 1 0 34500 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_365
timestamp 1644511149
transform 1 0 34684 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_377
timestamp 1644511149
transform 1 0 35788 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_389
timestamp 1644511149
transform 1 0 36892 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_401
timestamp 1644511149
transform 1 0 37996 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_413
timestamp 1644511149
transform 1 0 39100 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_419
timestamp 1644511149
transform 1 0 39652 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_421
timestamp 1644511149
transform 1 0 39836 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_433
timestamp 1644511149
transform 1 0 40940 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_445
timestamp 1644511149
transform 1 0 42044 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_457
timestamp 1644511149
transform 1 0 43148 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_469
timestamp 1644511149
transform 1 0 44252 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_475
timestamp 1644511149
transform 1 0 44804 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_477
timestamp 1644511149
transform 1 0 44988 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_489
timestamp 1644511149
transform 1 0 46092 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_501
timestamp 1644511149
transform 1 0 47196 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_513
timestamp 1644511149
transform 1 0 48300 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_525
timestamp 1644511149
transform 1 0 49404 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_531
timestamp 1644511149
transform 1 0 49956 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_533
timestamp 1644511149
transform 1 0 50140 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_545
timestamp 1644511149
transform 1 0 51244 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_557
timestamp 1644511149
transform 1 0 52348 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_569
timestamp 1644511149
transform 1 0 53452 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_581
timestamp 1644511149
transform 1 0 54556 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_587
timestamp 1644511149
transform 1 0 55108 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_589
timestamp 1644511149
transform 1 0 55292 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_601
timestamp 1644511149
transform 1 0 56396 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_609
timestamp 1644511149
transform 1 0 57132 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_613
timestamp 1644511149
transform 1 0 57500 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_3
timestamp 1644511149
transform 1 0 1380 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_15
timestamp 1644511149
transform 1 0 2484 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_27
timestamp 1644511149
transform 1 0 3588 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_39
timestamp 1644511149
transform 1 0 4692 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_51
timestamp 1644511149
transform 1 0 5796 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_55
timestamp 1644511149
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_57
timestamp 1644511149
transform 1 0 6348 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_69
timestamp 1644511149
transform 1 0 7452 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_81
timestamp 1644511149
transform 1 0 8556 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_93
timestamp 1644511149
transform 1 0 9660 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_105
timestamp 1644511149
transform 1 0 10764 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_111
timestamp 1644511149
transform 1 0 11316 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_113
timestamp 1644511149
transform 1 0 11500 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_125
timestamp 1644511149
transform 1 0 12604 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_137
timestamp 1644511149
transform 1 0 13708 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_149
timestamp 1644511149
transform 1 0 14812 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_161
timestamp 1644511149
transform 1 0 15916 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_167
timestamp 1644511149
transform 1 0 16468 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_169
timestamp 1644511149
transform 1 0 16652 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_181
timestamp 1644511149
transform 1 0 17756 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_193
timestamp 1644511149
transform 1 0 18860 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_205
timestamp 1644511149
transform 1 0 19964 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_217
timestamp 1644511149
transform 1 0 21068 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_223
timestamp 1644511149
transform 1 0 21620 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_225
timestamp 1644511149
transform 1 0 21804 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_237
timestamp 1644511149
transform 1 0 22908 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_249
timestamp 1644511149
transform 1 0 24012 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_261
timestamp 1644511149
transform 1 0 25116 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_273
timestamp 1644511149
transform 1 0 26220 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_279
timestamp 1644511149
transform 1 0 26772 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_281
timestamp 1644511149
transform 1 0 26956 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_293
timestamp 1644511149
transform 1 0 28060 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_305
timestamp 1644511149
transform 1 0 29164 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_317
timestamp 1644511149
transform 1 0 30268 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_329
timestamp 1644511149
transform 1 0 31372 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_335
timestamp 1644511149
transform 1 0 31924 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_337
timestamp 1644511149
transform 1 0 32108 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_349
timestamp 1644511149
transform 1 0 33212 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_361
timestamp 1644511149
transform 1 0 34316 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_373
timestamp 1644511149
transform 1 0 35420 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_385
timestamp 1644511149
transform 1 0 36524 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_391
timestamp 1644511149
transform 1 0 37076 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_393
timestamp 1644511149
transform 1 0 37260 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_405
timestamp 1644511149
transform 1 0 38364 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_417
timestamp 1644511149
transform 1 0 39468 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_429
timestamp 1644511149
transform 1 0 40572 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_441
timestamp 1644511149
transform 1 0 41676 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_447
timestamp 1644511149
transform 1 0 42228 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_449
timestamp 1644511149
transform 1 0 42412 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_461
timestamp 1644511149
transform 1 0 43516 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_473
timestamp 1644511149
transform 1 0 44620 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_485
timestamp 1644511149
transform 1 0 45724 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_497
timestamp 1644511149
transform 1 0 46828 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_503
timestamp 1644511149
transform 1 0 47380 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_505
timestamp 1644511149
transform 1 0 47564 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_517
timestamp 1644511149
transform 1 0 48668 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_529
timestamp 1644511149
transform 1 0 49772 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_541
timestamp 1644511149
transform 1 0 50876 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_553
timestamp 1644511149
transform 1 0 51980 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_559
timestamp 1644511149
transform 1 0 52532 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_561
timestamp 1644511149
transform 1 0 52716 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_573
timestamp 1644511149
transform 1 0 53820 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_585
timestamp 1644511149
transform 1 0 54924 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_597
timestamp 1644511149
transform 1 0 56028 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_609
timestamp 1644511149
transform 1 0 57132 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_615
timestamp 1644511149
transform 1 0 57684 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_617
timestamp 1644511149
transform 1 0 57868 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_20_3
timestamp 1644511149
transform 1 0 1380 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_15
timestamp 1644511149
transform 1 0 2484 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_27
timestamp 1644511149
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_29
timestamp 1644511149
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_41
timestamp 1644511149
transform 1 0 4876 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_53
timestamp 1644511149
transform 1 0 5980 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_65
timestamp 1644511149
transform 1 0 7084 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_77
timestamp 1644511149
transform 1 0 8188 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_83
timestamp 1644511149
transform 1 0 8740 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_85
timestamp 1644511149
transform 1 0 8924 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_97
timestamp 1644511149
transform 1 0 10028 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_109
timestamp 1644511149
transform 1 0 11132 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_121
timestamp 1644511149
transform 1 0 12236 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_133
timestamp 1644511149
transform 1 0 13340 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_139
timestamp 1644511149
transform 1 0 13892 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_141
timestamp 1644511149
transform 1 0 14076 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_153
timestamp 1644511149
transform 1 0 15180 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_165
timestamp 1644511149
transform 1 0 16284 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_177
timestamp 1644511149
transform 1 0 17388 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_189
timestamp 1644511149
transform 1 0 18492 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_195
timestamp 1644511149
transform 1 0 19044 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_197
timestamp 1644511149
transform 1 0 19228 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_209
timestamp 1644511149
transform 1 0 20332 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_221
timestamp 1644511149
transform 1 0 21436 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_233
timestamp 1644511149
transform 1 0 22540 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_245
timestamp 1644511149
transform 1 0 23644 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_251
timestamp 1644511149
transform 1 0 24196 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_253
timestamp 1644511149
transform 1 0 24380 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_265
timestamp 1644511149
transform 1 0 25484 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_277
timestamp 1644511149
transform 1 0 26588 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_289
timestamp 1644511149
transform 1 0 27692 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_301
timestamp 1644511149
transform 1 0 28796 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_307
timestamp 1644511149
transform 1 0 29348 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_309
timestamp 1644511149
transform 1 0 29532 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_321
timestamp 1644511149
transform 1 0 30636 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_333
timestamp 1644511149
transform 1 0 31740 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_345
timestamp 1644511149
transform 1 0 32844 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_357
timestamp 1644511149
transform 1 0 33948 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_363
timestamp 1644511149
transform 1 0 34500 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_365
timestamp 1644511149
transform 1 0 34684 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_377
timestamp 1644511149
transform 1 0 35788 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_389
timestamp 1644511149
transform 1 0 36892 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_401
timestamp 1644511149
transform 1 0 37996 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_413
timestamp 1644511149
transform 1 0 39100 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_419
timestamp 1644511149
transform 1 0 39652 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_421
timestamp 1644511149
transform 1 0 39836 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_433
timestamp 1644511149
transform 1 0 40940 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_445
timestamp 1644511149
transform 1 0 42044 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_457
timestamp 1644511149
transform 1 0 43148 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_469
timestamp 1644511149
transform 1 0 44252 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_475
timestamp 1644511149
transform 1 0 44804 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_477
timestamp 1644511149
transform 1 0 44988 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_489
timestamp 1644511149
transform 1 0 46092 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_501
timestamp 1644511149
transform 1 0 47196 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_513
timestamp 1644511149
transform 1 0 48300 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_525
timestamp 1644511149
transform 1 0 49404 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_531
timestamp 1644511149
transform 1 0 49956 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_533
timestamp 1644511149
transform 1 0 50140 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_545
timestamp 1644511149
transform 1 0 51244 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_557
timestamp 1644511149
transform 1 0 52348 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_569
timestamp 1644511149
transform 1 0 53452 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_581
timestamp 1644511149
transform 1 0 54556 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_587
timestamp 1644511149
transform 1 0 55108 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_589
timestamp 1644511149
transform 1 0 55292 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_601
timestamp 1644511149
transform 1 0 56396 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_613
timestamp 1644511149
transform 1 0 57500 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_3
timestamp 1644511149
transform 1 0 1380 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_15
timestamp 1644511149
transform 1 0 2484 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_27
timestamp 1644511149
transform 1 0 3588 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_39
timestamp 1644511149
transform 1 0 4692 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_51
timestamp 1644511149
transform 1 0 5796 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_55
timestamp 1644511149
transform 1 0 6164 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_57
timestamp 1644511149
transform 1 0 6348 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_69
timestamp 1644511149
transform 1 0 7452 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_81
timestamp 1644511149
transform 1 0 8556 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_93
timestamp 1644511149
transform 1 0 9660 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_105
timestamp 1644511149
transform 1 0 10764 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_111
timestamp 1644511149
transform 1 0 11316 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_113
timestamp 1644511149
transform 1 0 11500 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_125
timestamp 1644511149
transform 1 0 12604 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_137
timestamp 1644511149
transform 1 0 13708 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_149
timestamp 1644511149
transform 1 0 14812 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_161
timestamp 1644511149
transform 1 0 15916 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_167
timestamp 1644511149
transform 1 0 16468 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_169
timestamp 1644511149
transform 1 0 16652 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_181
timestamp 1644511149
transform 1 0 17756 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_193
timestamp 1644511149
transform 1 0 18860 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_205
timestamp 1644511149
transform 1 0 19964 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_217
timestamp 1644511149
transform 1 0 21068 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_223
timestamp 1644511149
transform 1 0 21620 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_225
timestamp 1644511149
transform 1 0 21804 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_237
timestamp 1644511149
transform 1 0 22908 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_249
timestamp 1644511149
transform 1 0 24012 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_261
timestamp 1644511149
transform 1 0 25116 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_273
timestamp 1644511149
transform 1 0 26220 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_279
timestamp 1644511149
transform 1 0 26772 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_281
timestamp 1644511149
transform 1 0 26956 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_293
timestamp 1644511149
transform 1 0 28060 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_305
timestamp 1644511149
transform 1 0 29164 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_317
timestamp 1644511149
transform 1 0 30268 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_329
timestamp 1644511149
transform 1 0 31372 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_335
timestamp 1644511149
transform 1 0 31924 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_337
timestamp 1644511149
transform 1 0 32108 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_349
timestamp 1644511149
transform 1 0 33212 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_361
timestamp 1644511149
transform 1 0 34316 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_373
timestamp 1644511149
transform 1 0 35420 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_385
timestamp 1644511149
transform 1 0 36524 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_391
timestamp 1644511149
transform 1 0 37076 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_393
timestamp 1644511149
transform 1 0 37260 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_405
timestamp 1644511149
transform 1 0 38364 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_417
timestamp 1644511149
transform 1 0 39468 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_429
timestamp 1644511149
transform 1 0 40572 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_441
timestamp 1644511149
transform 1 0 41676 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_447
timestamp 1644511149
transform 1 0 42228 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_449
timestamp 1644511149
transform 1 0 42412 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_461
timestamp 1644511149
transform 1 0 43516 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_473
timestamp 1644511149
transform 1 0 44620 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_485
timestamp 1644511149
transform 1 0 45724 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_497
timestamp 1644511149
transform 1 0 46828 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_503
timestamp 1644511149
transform 1 0 47380 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_505
timestamp 1644511149
transform 1 0 47564 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_517
timestamp 1644511149
transform 1 0 48668 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_529
timestamp 1644511149
transform 1 0 49772 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_541
timestamp 1644511149
transform 1 0 50876 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_553
timestamp 1644511149
transform 1 0 51980 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_559
timestamp 1644511149
transform 1 0 52532 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_561
timestamp 1644511149
transform 1 0 52716 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_573
timestamp 1644511149
transform 1 0 53820 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_585
timestamp 1644511149
transform 1 0 54924 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_597
timestamp 1644511149
transform 1 0 56028 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_609
timestamp 1644511149
transform 1 0 57132 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_615
timestamp 1644511149
transform 1 0 57684 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_617
timestamp 1644511149
transform 1 0 57868 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_22_3
timestamp 1644511149
transform 1 0 1380 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_15
timestamp 1644511149
transform 1 0 2484 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_27
timestamp 1644511149
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_29
timestamp 1644511149
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_41
timestamp 1644511149
transform 1 0 4876 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_53
timestamp 1644511149
transform 1 0 5980 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_65
timestamp 1644511149
transform 1 0 7084 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_77
timestamp 1644511149
transform 1 0 8188 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_83
timestamp 1644511149
transform 1 0 8740 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_85
timestamp 1644511149
transform 1 0 8924 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_97
timestamp 1644511149
transform 1 0 10028 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_109
timestamp 1644511149
transform 1 0 11132 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_121
timestamp 1644511149
transform 1 0 12236 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_133
timestamp 1644511149
transform 1 0 13340 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_139
timestamp 1644511149
transform 1 0 13892 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_141
timestamp 1644511149
transform 1 0 14076 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_153
timestamp 1644511149
transform 1 0 15180 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_165
timestamp 1644511149
transform 1 0 16284 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_177
timestamp 1644511149
transform 1 0 17388 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_189
timestamp 1644511149
transform 1 0 18492 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_195
timestamp 1644511149
transform 1 0 19044 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_197
timestamp 1644511149
transform 1 0 19228 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_209
timestamp 1644511149
transform 1 0 20332 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_221
timestamp 1644511149
transform 1 0 21436 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_233
timestamp 1644511149
transform 1 0 22540 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_245
timestamp 1644511149
transform 1 0 23644 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_251
timestamp 1644511149
transform 1 0 24196 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_253
timestamp 1644511149
transform 1 0 24380 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_265
timestamp 1644511149
transform 1 0 25484 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_277
timestamp 1644511149
transform 1 0 26588 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_289
timestamp 1644511149
transform 1 0 27692 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_301
timestamp 1644511149
transform 1 0 28796 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_307
timestamp 1644511149
transform 1 0 29348 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_309
timestamp 1644511149
transform 1 0 29532 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_321
timestamp 1644511149
transform 1 0 30636 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_333
timestamp 1644511149
transform 1 0 31740 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_345
timestamp 1644511149
transform 1 0 32844 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_357
timestamp 1644511149
transform 1 0 33948 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_363
timestamp 1644511149
transform 1 0 34500 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_365
timestamp 1644511149
transform 1 0 34684 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_377
timestamp 1644511149
transform 1 0 35788 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_389
timestamp 1644511149
transform 1 0 36892 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_401
timestamp 1644511149
transform 1 0 37996 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_413
timestamp 1644511149
transform 1 0 39100 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_419
timestamp 1644511149
transform 1 0 39652 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_421
timestamp 1644511149
transform 1 0 39836 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_433
timestamp 1644511149
transform 1 0 40940 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_445
timestamp 1644511149
transform 1 0 42044 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_457
timestamp 1644511149
transform 1 0 43148 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_469
timestamp 1644511149
transform 1 0 44252 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_475
timestamp 1644511149
transform 1 0 44804 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_477
timestamp 1644511149
transform 1 0 44988 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_489
timestamp 1644511149
transform 1 0 46092 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_501
timestamp 1644511149
transform 1 0 47196 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_513
timestamp 1644511149
transform 1 0 48300 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_525
timestamp 1644511149
transform 1 0 49404 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_531
timestamp 1644511149
transform 1 0 49956 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_533
timestamp 1644511149
transform 1 0 50140 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_545
timestamp 1644511149
transform 1 0 51244 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_557
timestamp 1644511149
transform 1 0 52348 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_569
timestamp 1644511149
transform 1 0 53452 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_581
timestamp 1644511149
transform 1 0 54556 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_587
timestamp 1644511149
transform 1 0 55108 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_589
timestamp 1644511149
transform 1 0 55292 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_601
timestamp 1644511149
transform 1 0 56396 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_613
timestamp 1644511149
transform 1 0 57500 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_3
timestamp 1644511149
transform 1 0 1380 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_15
timestamp 1644511149
transform 1 0 2484 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_27
timestamp 1644511149
transform 1 0 3588 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_39
timestamp 1644511149
transform 1 0 4692 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_51
timestamp 1644511149
transform 1 0 5796 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_55
timestamp 1644511149
transform 1 0 6164 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_57
timestamp 1644511149
transform 1 0 6348 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_69
timestamp 1644511149
transform 1 0 7452 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_81
timestamp 1644511149
transform 1 0 8556 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_93
timestamp 1644511149
transform 1 0 9660 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_105
timestamp 1644511149
transform 1 0 10764 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_111
timestamp 1644511149
transform 1 0 11316 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_113
timestamp 1644511149
transform 1 0 11500 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_125
timestamp 1644511149
transform 1 0 12604 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_137
timestamp 1644511149
transform 1 0 13708 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_149
timestamp 1644511149
transform 1 0 14812 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_161
timestamp 1644511149
transform 1 0 15916 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_167
timestamp 1644511149
transform 1 0 16468 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_169
timestamp 1644511149
transform 1 0 16652 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_181
timestamp 1644511149
transform 1 0 17756 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_193
timestamp 1644511149
transform 1 0 18860 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_205
timestamp 1644511149
transform 1 0 19964 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_217
timestamp 1644511149
transform 1 0 21068 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_223
timestamp 1644511149
transform 1 0 21620 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_225
timestamp 1644511149
transform 1 0 21804 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_237
timestamp 1644511149
transform 1 0 22908 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_249
timestamp 1644511149
transform 1 0 24012 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_261
timestamp 1644511149
transform 1 0 25116 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_273
timestamp 1644511149
transform 1 0 26220 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_279
timestamp 1644511149
transform 1 0 26772 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_281
timestamp 1644511149
transform 1 0 26956 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_293
timestamp 1644511149
transform 1 0 28060 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_305
timestamp 1644511149
transform 1 0 29164 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_317
timestamp 1644511149
transform 1 0 30268 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_329
timestamp 1644511149
transform 1 0 31372 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_335
timestamp 1644511149
transform 1 0 31924 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_337
timestamp 1644511149
transform 1 0 32108 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_349
timestamp 1644511149
transform 1 0 33212 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_361
timestamp 1644511149
transform 1 0 34316 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_373
timestamp 1644511149
transform 1 0 35420 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_385
timestamp 1644511149
transform 1 0 36524 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_391
timestamp 1644511149
transform 1 0 37076 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_393
timestamp 1644511149
transform 1 0 37260 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_405
timestamp 1644511149
transform 1 0 38364 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_417
timestamp 1644511149
transform 1 0 39468 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_429
timestamp 1644511149
transform 1 0 40572 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_441
timestamp 1644511149
transform 1 0 41676 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_447
timestamp 1644511149
transform 1 0 42228 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_449
timestamp 1644511149
transform 1 0 42412 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_461
timestamp 1644511149
transform 1 0 43516 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_473
timestamp 1644511149
transform 1 0 44620 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_485
timestamp 1644511149
transform 1 0 45724 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_497
timestamp 1644511149
transform 1 0 46828 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_503
timestamp 1644511149
transform 1 0 47380 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_505
timestamp 1644511149
transform 1 0 47564 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_517
timestamp 1644511149
transform 1 0 48668 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_529
timestamp 1644511149
transform 1 0 49772 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_541
timestamp 1644511149
transform 1 0 50876 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_553
timestamp 1644511149
transform 1 0 51980 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_559
timestamp 1644511149
transform 1 0 52532 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_561
timestamp 1644511149
transform 1 0 52716 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_573
timestamp 1644511149
transform 1 0 53820 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_585
timestamp 1644511149
transform 1 0 54924 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_597
timestamp 1644511149
transform 1 0 56028 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_609
timestamp 1644511149
transform 1 0 57132 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_615
timestamp 1644511149
transform 1 0 57684 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_617
timestamp 1644511149
transform 1 0 57868 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_24_3
timestamp 1644511149
transform 1 0 1380 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_15
timestamp 1644511149
transform 1 0 2484 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_27
timestamp 1644511149
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_29
timestamp 1644511149
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_41
timestamp 1644511149
transform 1 0 4876 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_53
timestamp 1644511149
transform 1 0 5980 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_65
timestamp 1644511149
transform 1 0 7084 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_77
timestamp 1644511149
transform 1 0 8188 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_83
timestamp 1644511149
transform 1 0 8740 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_85
timestamp 1644511149
transform 1 0 8924 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_97
timestamp 1644511149
transform 1 0 10028 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_109
timestamp 1644511149
transform 1 0 11132 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_121
timestamp 1644511149
transform 1 0 12236 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_133
timestamp 1644511149
transform 1 0 13340 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_139
timestamp 1644511149
transform 1 0 13892 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_141
timestamp 1644511149
transform 1 0 14076 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_153
timestamp 1644511149
transform 1 0 15180 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_165
timestamp 1644511149
transform 1 0 16284 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_177
timestamp 1644511149
transform 1 0 17388 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_189
timestamp 1644511149
transform 1 0 18492 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_195
timestamp 1644511149
transform 1 0 19044 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_197
timestamp 1644511149
transform 1 0 19228 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_209
timestamp 1644511149
transform 1 0 20332 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_221
timestamp 1644511149
transform 1 0 21436 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_233
timestamp 1644511149
transform 1 0 22540 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_245
timestamp 1644511149
transform 1 0 23644 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_251
timestamp 1644511149
transform 1 0 24196 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_253
timestamp 1644511149
transform 1 0 24380 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_265
timestamp 1644511149
transform 1 0 25484 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_277
timestamp 1644511149
transform 1 0 26588 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_289
timestamp 1644511149
transform 1 0 27692 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_301
timestamp 1644511149
transform 1 0 28796 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_307
timestamp 1644511149
transform 1 0 29348 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_309
timestamp 1644511149
transform 1 0 29532 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_321
timestamp 1644511149
transform 1 0 30636 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_333
timestamp 1644511149
transform 1 0 31740 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_345
timestamp 1644511149
transform 1 0 32844 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_357
timestamp 1644511149
transform 1 0 33948 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_363
timestamp 1644511149
transform 1 0 34500 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_365
timestamp 1644511149
transform 1 0 34684 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_377
timestamp 1644511149
transform 1 0 35788 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_389
timestamp 1644511149
transform 1 0 36892 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_401
timestamp 1644511149
transform 1 0 37996 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_413
timestamp 1644511149
transform 1 0 39100 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_419
timestamp 1644511149
transform 1 0 39652 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_421
timestamp 1644511149
transform 1 0 39836 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_433
timestamp 1644511149
transform 1 0 40940 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_445
timestamp 1644511149
transform 1 0 42044 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_457
timestamp 1644511149
transform 1 0 43148 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_469
timestamp 1644511149
transform 1 0 44252 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_475
timestamp 1644511149
transform 1 0 44804 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_477
timestamp 1644511149
transform 1 0 44988 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_489
timestamp 1644511149
transform 1 0 46092 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_501
timestamp 1644511149
transform 1 0 47196 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_513
timestamp 1644511149
transform 1 0 48300 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_525
timestamp 1644511149
transform 1 0 49404 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_531
timestamp 1644511149
transform 1 0 49956 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_533
timestamp 1644511149
transform 1 0 50140 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_545
timestamp 1644511149
transform 1 0 51244 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_557
timestamp 1644511149
transform 1 0 52348 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_569
timestamp 1644511149
transform 1 0 53452 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_581
timestamp 1644511149
transform 1 0 54556 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_587
timestamp 1644511149
transform 1 0 55108 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_589
timestamp 1644511149
transform 1 0 55292 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_601
timestamp 1644511149
transform 1 0 56396 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_613
timestamp 1644511149
transform 1 0 57500 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_3
timestamp 1644511149
transform 1 0 1380 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_15
timestamp 1644511149
transform 1 0 2484 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_27
timestamp 1644511149
transform 1 0 3588 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_39
timestamp 1644511149
transform 1 0 4692 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_51
timestamp 1644511149
transform 1 0 5796 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_55
timestamp 1644511149
transform 1 0 6164 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_57
timestamp 1644511149
transform 1 0 6348 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_69
timestamp 1644511149
transform 1 0 7452 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_81
timestamp 1644511149
transform 1 0 8556 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_93
timestamp 1644511149
transform 1 0 9660 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_105
timestamp 1644511149
transform 1 0 10764 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_111
timestamp 1644511149
transform 1 0 11316 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_113
timestamp 1644511149
transform 1 0 11500 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_125
timestamp 1644511149
transform 1 0 12604 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_137
timestamp 1644511149
transform 1 0 13708 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_149
timestamp 1644511149
transform 1 0 14812 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_161
timestamp 1644511149
transform 1 0 15916 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_167
timestamp 1644511149
transform 1 0 16468 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_169
timestamp 1644511149
transform 1 0 16652 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_181
timestamp 1644511149
transform 1 0 17756 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_193
timestamp 1644511149
transform 1 0 18860 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_205
timestamp 1644511149
transform 1 0 19964 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_217
timestamp 1644511149
transform 1 0 21068 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_223
timestamp 1644511149
transform 1 0 21620 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_225
timestamp 1644511149
transform 1 0 21804 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_237
timestamp 1644511149
transform 1 0 22908 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_249
timestamp 1644511149
transform 1 0 24012 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_261
timestamp 1644511149
transform 1 0 25116 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_273
timestamp 1644511149
transform 1 0 26220 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_279
timestamp 1644511149
transform 1 0 26772 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_281
timestamp 1644511149
transform 1 0 26956 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_293
timestamp 1644511149
transform 1 0 28060 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_305
timestamp 1644511149
transform 1 0 29164 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_317
timestamp 1644511149
transform 1 0 30268 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_329
timestamp 1644511149
transform 1 0 31372 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_335
timestamp 1644511149
transform 1 0 31924 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_337
timestamp 1644511149
transform 1 0 32108 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_349
timestamp 1644511149
transform 1 0 33212 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_361
timestamp 1644511149
transform 1 0 34316 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_373
timestamp 1644511149
transform 1 0 35420 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_385
timestamp 1644511149
transform 1 0 36524 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_391
timestamp 1644511149
transform 1 0 37076 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_393
timestamp 1644511149
transform 1 0 37260 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_405
timestamp 1644511149
transform 1 0 38364 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_417
timestamp 1644511149
transform 1 0 39468 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_429
timestamp 1644511149
transform 1 0 40572 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_441
timestamp 1644511149
transform 1 0 41676 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_447
timestamp 1644511149
transform 1 0 42228 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_449
timestamp 1644511149
transform 1 0 42412 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_461
timestamp 1644511149
transform 1 0 43516 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_473
timestamp 1644511149
transform 1 0 44620 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_485
timestamp 1644511149
transform 1 0 45724 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_497
timestamp 1644511149
transform 1 0 46828 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_503
timestamp 1644511149
transform 1 0 47380 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_505
timestamp 1644511149
transform 1 0 47564 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_517
timestamp 1644511149
transform 1 0 48668 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_529
timestamp 1644511149
transform 1 0 49772 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_541
timestamp 1644511149
transform 1 0 50876 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_553
timestamp 1644511149
transform 1 0 51980 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_559
timestamp 1644511149
transform 1 0 52532 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_561
timestamp 1644511149
transform 1 0 52716 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_573
timestamp 1644511149
transform 1 0 53820 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_585
timestamp 1644511149
transform 1 0 54924 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_597
timestamp 1644511149
transform 1 0 56028 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_609
timestamp 1644511149
transform 1 0 57132 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_615
timestamp 1644511149
transform 1 0 57684 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_617
timestamp 1644511149
transform 1 0 57868 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_26_3
timestamp 1644511149
transform 1 0 1380 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_15
timestamp 1644511149
transform 1 0 2484 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_27
timestamp 1644511149
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_29
timestamp 1644511149
transform 1 0 3772 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_41
timestamp 1644511149
transform 1 0 4876 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_53
timestamp 1644511149
transform 1 0 5980 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_65
timestamp 1644511149
transform 1 0 7084 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_77
timestamp 1644511149
transform 1 0 8188 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_83
timestamp 1644511149
transform 1 0 8740 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_85
timestamp 1644511149
transform 1 0 8924 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_97
timestamp 1644511149
transform 1 0 10028 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_109
timestamp 1644511149
transform 1 0 11132 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_121
timestamp 1644511149
transform 1 0 12236 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_133
timestamp 1644511149
transform 1 0 13340 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_139
timestamp 1644511149
transform 1 0 13892 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_141
timestamp 1644511149
transform 1 0 14076 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_153
timestamp 1644511149
transform 1 0 15180 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_165
timestamp 1644511149
transform 1 0 16284 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_177
timestamp 1644511149
transform 1 0 17388 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_189
timestamp 1644511149
transform 1 0 18492 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_195
timestamp 1644511149
transform 1 0 19044 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_197
timestamp 1644511149
transform 1 0 19228 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_209
timestamp 1644511149
transform 1 0 20332 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_221
timestamp 1644511149
transform 1 0 21436 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_233
timestamp 1644511149
transform 1 0 22540 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_245
timestamp 1644511149
transform 1 0 23644 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_251
timestamp 1644511149
transform 1 0 24196 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_253
timestamp 1644511149
transform 1 0 24380 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_265
timestamp 1644511149
transform 1 0 25484 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_277
timestamp 1644511149
transform 1 0 26588 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_289
timestamp 1644511149
transform 1 0 27692 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_301
timestamp 1644511149
transform 1 0 28796 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_307
timestamp 1644511149
transform 1 0 29348 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_309
timestamp 1644511149
transform 1 0 29532 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_321
timestamp 1644511149
transform 1 0 30636 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_333
timestamp 1644511149
transform 1 0 31740 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_345
timestamp 1644511149
transform 1 0 32844 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_357
timestamp 1644511149
transform 1 0 33948 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_363
timestamp 1644511149
transform 1 0 34500 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_365
timestamp 1644511149
transform 1 0 34684 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_377
timestamp 1644511149
transform 1 0 35788 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_389
timestamp 1644511149
transform 1 0 36892 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_401
timestamp 1644511149
transform 1 0 37996 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_413
timestamp 1644511149
transform 1 0 39100 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_419
timestamp 1644511149
transform 1 0 39652 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_421
timestamp 1644511149
transform 1 0 39836 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_433
timestamp 1644511149
transform 1 0 40940 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_445
timestamp 1644511149
transform 1 0 42044 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_457
timestamp 1644511149
transform 1 0 43148 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_469
timestamp 1644511149
transform 1 0 44252 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_475
timestamp 1644511149
transform 1 0 44804 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_477
timestamp 1644511149
transform 1 0 44988 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_489
timestamp 1644511149
transform 1 0 46092 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_501
timestamp 1644511149
transform 1 0 47196 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_513
timestamp 1644511149
transform 1 0 48300 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_525
timestamp 1644511149
transform 1 0 49404 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_531
timestamp 1644511149
transform 1 0 49956 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_533
timestamp 1644511149
transform 1 0 50140 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_545
timestamp 1644511149
transform 1 0 51244 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_557
timestamp 1644511149
transform 1 0 52348 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_569
timestamp 1644511149
transform 1 0 53452 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_581
timestamp 1644511149
transform 1 0 54556 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_587
timestamp 1644511149
transform 1 0 55108 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_589
timestamp 1644511149
transform 1 0 55292 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_601
timestamp 1644511149
transform 1 0 56396 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_613
timestamp 1644511149
transform 1 0 57500 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_3
timestamp 1644511149
transform 1 0 1380 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_15
timestamp 1644511149
transform 1 0 2484 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_27
timestamp 1644511149
transform 1 0 3588 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_39
timestamp 1644511149
transform 1 0 4692 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_51
timestamp 1644511149
transform 1 0 5796 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_55
timestamp 1644511149
transform 1 0 6164 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_57
timestamp 1644511149
transform 1 0 6348 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_69
timestamp 1644511149
transform 1 0 7452 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_81
timestamp 1644511149
transform 1 0 8556 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_93
timestamp 1644511149
transform 1 0 9660 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_105
timestamp 1644511149
transform 1 0 10764 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_111
timestamp 1644511149
transform 1 0 11316 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_113
timestamp 1644511149
transform 1 0 11500 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_125
timestamp 1644511149
transform 1 0 12604 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_137
timestamp 1644511149
transform 1 0 13708 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_149
timestamp 1644511149
transform 1 0 14812 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_161
timestamp 1644511149
transform 1 0 15916 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_167
timestamp 1644511149
transform 1 0 16468 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_169
timestamp 1644511149
transform 1 0 16652 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_181
timestamp 1644511149
transform 1 0 17756 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_193
timestamp 1644511149
transform 1 0 18860 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_205
timestamp 1644511149
transform 1 0 19964 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_217
timestamp 1644511149
transform 1 0 21068 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_223
timestamp 1644511149
transform 1 0 21620 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_225
timestamp 1644511149
transform 1 0 21804 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_237
timestamp 1644511149
transform 1 0 22908 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_249
timestamp 1644511149
transform 1 0 24012 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_261
timestamp 1644511149
transform 1 0 25116 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_273
timestamp 1644511149
transform 1 0 26220 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_279
timestamp 1644511149
transform 1 0 26772 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_281
timestamp 1644511149
transform 1 0 26956 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_293
timestamp 1644511149
transform 1 0 28060 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_305
timestamp 1644511149
transform 1 0 29164 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_317
timestamp 1644511149
transform 1 0 30268 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_329
timestamp 1644511149
transform 1 0 31372 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_335
timestamp 1644511149
transform 1 0 31924 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_337
timestamp 1644511149
transform 1 0 32108 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_349
timestamp 1644511149
transform 1 0 33212 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_361
timestamp 1644511149
transform 1 0 34316 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_373
timestamp 1644511149
transform 1 0 35420 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_385
timestamp 1644511149
transform 1 0 36524 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_391
timestamp 1644511149
transform 1 0 37076 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_393
timestamp 1644511149
transform 1 0 37260 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_405
timestamp 1644511149
transform 1 0 38364 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_417
timestamp 1644511149
transform 1 0 39468 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_429
timestamp 1644511149
transform 1 0 40572 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_441
timestamp 1644511149
transform 1 0 41676 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_447
timestamp 1644511149
transform 1 0 42228 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_449
timestamp 1644511149
transform 1 0 42412 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_461
timestamp 1644511149
transform 1 0 43516 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_473
timestamp 1644511149
transform 1 0 44620 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_485
timestamp 1644511149
transform 1 0 45724 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_497
timestamp 1644511149
transform 1 0 46828 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_503
timestamp 1644511149
transform 1 0 47380 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_505
timestamp 1644511149
transform 1 0 47564 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_517
timestamp 1644511149
transform 1 0 48668 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_529
timestamp 1644511149
transform 1 0 49772 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_541
timestamp 1644511149
transform 1 0 50876 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_553
timestamp 1644511149
transform 1 0 51980 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_559
timestamp 1644511149
transform 1 0 52532 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_561
timestamp 1644511149
transform 1 0 52716 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_573
timestamp 1644511149
transform 1 0 53820 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_585
timestamp 1644511149
transform 1 0 54924 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_597
timestamp 1644511149
transform 1 0 56028 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_609
timestamp 1644511149
transform 1 0 57132 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_615
timestamp 1644511149
transform 1 0 57684 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_27_617
timestamp 1644511149
transform 1 0 57868 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_28_3
timestamp 1644511149
transform 1 0 1380 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_15
timestamp 1644511149
transform 1 0 2484 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_27
timestamp 1644511149
transform 1 0 3588 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_29
timestamp 1644511149
transform 1 0 3772 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_41
timestamp 1644511149
transform 1 0 4876 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_53
timestamp 1644511149
transform 1 0 5980 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_65
timestamp 1644511149
transform 1 0 7084 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_77
timestamp 1644511149
transform 1 0 8188 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_83
timestamp 1644511149
transform 1 0 8740 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_85
timestamp 1644511149
transform 1 0 8924 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_97
timestamp 1644511149
transform 1 0 10028 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_109
timestamp 1644511149
transform 1 0 11132 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_121
timestamp 1644511149
transform 1 0 12236 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_133
timestamp 1644511149
transform 1 0 13340 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_139
timestamp 1644511149
transform 1 0 13892 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_141
timestamp 1644511149
transform 1 0 14076 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_153
timestamp 1644511149
transform 1 0 15180 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_165
timestamp 1644511149
transform 1 0 16284 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_177
timestamp 1644511149
transform 1 0 17388 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_189
timestamp 1644511149
transform 1 0 18492 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_195
timestamp 1644511149
transform 1 0 19044 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_197
timestamp 1644511149
transform 1 0 19228 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_209
timestamp 1644511149
transform 1 0 20332 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_221
timestamp 1644511149
transform 1 0 21436 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_233
timestamp 1644511149
transform 1 0 22540 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_245
timestamp 1644511149
transform 1 0 23644 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_251
timestamp 1644511149
transform 1 0 24196 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_253
timestamp 1644511149
transform 1 0 24380 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_265
timestamp 1644511149
transform 1 0 25484 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_277
timestamp 1644511149
transform 1 0 26588 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_289
timestamp 1644511149
transform 1 0 27692 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_301
timestamp 1644511149
transform 1 0 28796 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_307
timestamp 1644511149
transform 1 0 29348 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_309
timestamp 1644511149
transform 1 0 29532 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_321
timestamp 1644511149
transform 1 0 30636 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_333
timestamp 1644511149
transform 1 0 31740 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_345
timestamp 1644511149
transform 1 0 32844 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_357
timestamp 1644511149
transform 1 0 33948 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_363
timestamp 1644511149
transform 1 0 34500 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_365
timestamp 1644511149
transform 1 0 34684 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_377
timestamp 1644511149
transform 1 0 35788 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_389
timestamp 1644511149
transform 1 0 36892 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_401
timestamp 1644511149
transform 1 0 37996 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_413
timestamp 1644511149
transform 1 0 39100 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_419
timestamp 1644511149
transform 1 0 39652 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_421
timestamp 1644511149
transform 1 0 39836 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_433
timestamp 1644511149
transform 1 0 40940 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_445
timestamp 1644511149
transform 1 0 42044 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_457
timestamp 1644511149
transform 1 0 43148 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_469
timestamp 1644511149
transform 1 0 44252 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_475
timestamp 1644511149
transform 1 0 44804 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_477
timestamp 1644511149
transform 1 0 44988 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_489
timestamp 1644511149
transform 1 0 46092 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_501
timestamp 1644511149
transform 1 0 47196 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_513
timestamp 1644511149
transform 1 0 48300 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_525
timestamp 1644511149
transform 1 0 49404 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_531
timestamp 1644511149
transform 1 0 49956 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_533
timestamp 1644511149
transform 1 0 50140 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_545
timestamp 1644511149
transform 1 0 51244 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_557
timestamp 1644511149
transform 1 0 52348 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_569
timestamp 1644511149
transform 1 0 53452 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_581
timestamp 1644511149
transform 1 0 54556 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_587
timestamp 1644511149
transform 1 0 55108 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_589
timestamp 1644511149
transform 1 0 55292 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_601
timestamp 1644511149
transform 1 0 56396 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_613
timestamp 1644511149
transform 1 0 57500 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_3
timestamp 1644511149
transform 1 0 1380 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_15
timestamp 1644511149
transform 1 0 2484 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_27
timestamp 1644511149
transform 1 0 3588 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_39
timestamp 1644511149
transform 1 0 4692 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_51
timestamp 1644511149
transform 1 0 5796 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_55
timestamp 1644511149
transform 1 0 6164 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_57
timestamp 1644511149
transform 1 0 6348 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_69
timestamp 1644511149
transform 1 0 7452 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_81
timestamp 1644511149
transform 1 0 8556 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_93
timestamp 1644511149
transform 1 0 9660 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_105
timestamp 1644511149
transform 1 0 10764 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_111
timestamp 1644511149
transform 1 0 11316 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_113
timestamp 1644511149
transform 1 0 11500 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_125
timestamp 1644511149
transform 1 0 12604 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_137
timestamp 1644511149
transform 1 0 13708 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_149
timestamp 1644511149
transform 1 0 14812 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_161
timestamp 1644511149
transform 1 0 15916 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_167
timestamp 1644511149
transform 1 0 16468 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_169
timestamp 1644511149
transform 1 0 16652 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_181
timestamp 1644511149
transform 1 0 17756 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_193
timestamp 1644511149
transform 1 0 18860 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_205
timestamp 1644511149
transform 1 0 19964 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_217
timestamp 1644511149
transform 1 0 21068 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_223
timestamp 1644511149
transform 1 0 21620 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_225
timestamp 1644511149
transform 1 0 21804 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_237
timestamp 1644511149
transform 1 0 22908 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_249
timestamp 1644511149
transform 1 0 24012 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_261
timestamp 1644511149
transform 1 0 25116 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_273
timestamp 1644511149
transform 1 0 26220 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_279
timestamp 1644511149
transform 1 0 26772 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_281
timestamp 1644511149
transform 1 0 26956 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_293
timestamp 1644511149
transform 1 0 28060 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_305
timestamp 1644511149
transform 1 0 29164 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_317
timestamp 1644511149
transform 1 0 30268 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_329
timestamp 1644511149
transform 1 0 31372 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_335
timestamp 1644511149
transform 1 0 31924 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_337
timestamp 1644511149
transform 1 0 32108 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_349
timestamp 1644511149
transform 1 0 33212 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_361
timestamp 1644511149
transform 1 0 34316 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_373
timestamp 1644511149
transform 1 0 35420 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_385
timestamp 1644511149
transform 1 0 36524 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_391
timestamp 1644511149
transform 1 0 37076 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_393
timestamp 1644511149
transform 1 0 37260 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_405
timestamp 1644511149
transform 1 0 38364 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_417
timestamp 1644511149
transform 1 0 39468 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_429
timestamp 1644511149
transform 1 0 40572 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_441
timestamp 1644511149
transform 1 0 41676 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_447
timestamp 1644511149
transform 1 0 42228 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_449
timestamp 1644511149
transform 1 0 42412 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_461
timestamp 1644511149
transform 1 0 43516 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_473
timestamp 1644511149
transform 1 0 44620 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_485
timestamp 1644511149
transform 1 0 45724 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_497
timestamp 1644511149
transform 1 0 46828 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_503
timestamp 1644511149
transform 1 0 47380 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_505
timestamp 1644511149
transform 1 0 47564 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_517
timestamp 1644511149
transform 1 0 48668 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_529
timestamp 1644511149
transform 1 0 49772 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_541
timestamp 1644511149
transform 1 0 50876 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_553
timestamp 1644511149
transform 1 0 51980 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_559
timestamp 1644511149
transform 1 0 52532 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_561
timestamp 1644511149
transform 1 0 52716 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_573
timestamp 1644511149
transform 1 0 53820 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_585
timestamp 1644511149
transform 1 0 54924 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_597
timestamp 1644511149
transform 1 0 56028 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_609
timestamp 1644511149
transform 1 0 57132 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_615
timestamp 1644511149
transform 1 0 57684 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_617
timestamp 1644511149
transform 1 0 57868 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_30_3
timestamp 1644511149
transform 1 0 1380 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_15
timestamp 1644511149
transform 1 0 2484 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_27
timestamp 1644511149
transform 1 0 3588 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_29
timestamp 1644511149
transform 1 0 3772 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_41
timestamp 1644511149
transform 1 0 4876 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_53
timestamp 1644511149
transform 1 0 5980 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_65
timestamp 1644511149
transform 1 0 7084 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_77
timestamp 1644511149
transform 1 0 8188 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_83
timestamp 1644511149
transform 1 0 8740 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_85
timestamp 1644511149
transform 1 0 8924 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_97
timestamp 1644511149
transform 1 0 10028 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_109
timestamp 1644511149
transform 1 0 11132 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_121
timestamp 1644511149
transform 1 0 12236 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_133
timestamp 1644511149
transform 1 0 13340 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_139
timestamp 1644511149
transform 1 0 13892 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_141
timestamp 1644511149
transform 1 0 14076 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_153
timestamp 1644511149
transform 1 0 15180 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_165
timestamp 1644511149
transform 1 0 16284 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_177
timestamp 1644511149
transform 1 0 17388 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_189
timestamp 1644511149
transform 1 0 18492 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_195
timestamp 1644511149
transform 1 0 19044 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_197
timestamp 1644511149
transform 1 0 19228 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_209
timestamp 1644511149
transform 1 0 20332 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_221
timestamp 1644511149
transform 1 0 21436 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_233
timestamp 1644511149
transform 1 0 22540 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_245
timestamp 1644511149
transform 1 0 23644 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_251
timestamp 1644511149
transform 1 0 24196 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_253
timestamp 1644511149
transform 1 0 24380 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_265
timestamp 1644511149
transform 1 0 25484 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_277
timestamp 1644511149
transform 1 0 26588 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_289
timestamp 1644511149
transform 1 0 27692 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_301
timestamp 1644511149
transform 1 0 28796 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_307
timestamp 1644511149
transform 1 0 29348 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_309
timestamp 1644511149
transform 1 0 29532 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_321
timestamp 1644511149
transform 1 0 30636 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_333
timestamp 1644511149
transform 1 0 31740 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_345
timestamp 1644511149
transform 1 0 32844 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_357
timestamp 1644511149
transform 1 0 33948 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_363
timestamp 1644511149
transform 1 0 34500 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_365
timestamp 1644511149
transform 1 0 34684 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_377
timestamp 1644511149
transform 1 0 35788 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_389
timestamp 1644511149
transform 1 0 36892 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_401
timestamp 1644511149
transform 1 0 37996 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_413
timestamp 1644511149
transform 1 0 39100 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_419
timestamp 1644511149
transform 1 0 39652 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_421
timestamp 1644511149
transform 1 0 39836 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_433
timestamp 1644511149
transform 1 0 40940 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_445
timestamp 1644511149
transform 1 0 42044 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_457
timestamp 1644511149
transform 1 0 43148 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_469
timestamp 1644511149
transform 1 0 44252 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_475
timestamp 1644511149
transform 1 0 44804 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_477
timestamp 1644511149
transform 1 0 44988 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_489
timestamp 1644511149
transform 1 0 46092 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_501
timestamp 1644511149
transform 1 0 47196 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_513
timestamp 1644511149
transform 1 0 48300 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_525
timestamp 1644511149
transform 1 0 49404 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_531
timestamp 1644511149
transform 1 0 49956 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_533
timestamp 1644511149
transform 1 0 50140 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_545
timestamp 1644511149
transform 1 0 51244 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_557
timestamp 1644511149
transform 1 0 52348 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_569
timestamp 1644511149
transform 1 0 53452 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_581
timestamp 1644511149
transform 1 0 54556 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_587
timestamp 1644511149
transform 1 0 55108 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_30_589
timestamp 1644511149
transform 1 0 55292 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_30_597
timestamp 1644511149
transform 1 0 56028 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_30_621
timestamp 1644511149
transform 1 0 58236 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_31_3
timestamp 1644511149
transform 1 0 1380 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_15
timestamp 1644511149
transform 1 0 2484 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_27
timestamp 1644511149
transform 1 0 3588 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_39
timestamp 1644511149
transform 1 0 4692 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_51
timestamp 1644511149
transform 1 0 5796 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_55
timestamp 1644511149
transform 1 0 6164 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_57
timestamp 1644511149
transform 1 0 6348 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_69
timestamp 1644511149
transform 1 0 7452 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_81
timestamp 1644511149
transform 1 0 8556 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_93
timestamp 1644511149
transform 1 0 9660 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_105
timestamp 1644511149
transform 1 0 10764 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_111
timestamp 1644511149
transform 1 0 11316 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_113
timestamp 1644511149
transform 1 0 11500 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_125
timestamp 1644511149
transform 1 0 12604 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_137
timestamp 1644511149
transform 1 0 13708 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_149
timestamp 1644511149
transform 1 0 14812 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_161
timestamp 1644511149
transform 1 0 15916 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_167
timestamp 1644511149
transform 1 0 16468 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_169
timestamp 1644511149
transform 1 0 16652 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_181
timestamp 1644511149
transform 1 0 17756 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_193
timestamp 1644511149
transform 1 0 18860 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_205
timestamp 1644511149
transform 1 0 19964 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_217
timestamp 1644511149
transform 1 0 21068 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_223
timestamp 1644511149
transform 1 0 21620 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_225
timestamp 1644511149
transform 1 0 21804 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_237
timestamp 1644511149
transform 1 0 22908 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_249
timestamp 1644511149
transform 1 0 24012 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_261
timestamp 1644511149
transform 1 0 25116 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_273
timestamp 1644511149
transform 1 0 26220 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_279
timestamp 1644511149
transform 1 0 26772 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_281
timestamp 1644511149
transform 1 0 26956 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_293
timestamp 1644511149
transform 1 0 28060 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_305
timestamp 1644511149
transform 1 0 29164 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_317
timestamp 1644511149
transform 1 0 30268 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_329
timestamp 1644511149
transform 1 0 31372 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_335
timestamp 1644511149
transform 1 0 31924 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_337
timestamp 1644511149
transform 1 0 32108 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_349
timestamp 1644511149
transform 1 0 33212 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_361
timestamp 1644511149
transform 1 0 34316 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_373
timestamp 1644511149
transform 1 0 35420 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_385
timestamp 1644511149
transform 1 0 36524 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_391
timestamp 1644511149
transform 1 0 37076 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_393
timestamp 1644511149
transform 1 0 37260 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_405
timestamp 1644511149
transform 1 0 38364 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_417
timestamp 1644511149
transform 1 0 39468 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_429
timestamp 1644511149
transform 1 0 40572 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_441
timestamp 1644511149
transform 1 0 41676 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_447
timestamp 1644511149
transform 1 0 42228 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_449
timestamp 1644511149
transform 1 0 42412 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_461
timestamp 1644511149
transform 1 0 43516 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_473
timestamp 1644511149
transform 1 0 44620 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_485
timestamp 1644511149
transform 1 0 45724 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_497
timestamp 1644511149
transform 1 0 46828 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_503
timestamp 1644511149
transform 1 0 47380 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_505
timestamp 1644511149
transform 1 0 47564 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_517
timestamp 1644511149
transform 1 0 48668 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_529
timestamp 1644511149
transform 1 0 49772 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_541
timestamp 1644511149
transform 1 0 50876 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_553
timestamp 1644511149
transform 1 0 51980 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_559
timestamp 1644511149
transform 1 0 52532 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_561
timestamp 1644511149
transform 1 0 52716 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_573
timestamp 1644511149
transform 1 0 53820 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_585
timestamp 1644511149
transform 1 0 54924 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_31_597
timestamp 1644511149
transform 1 0 56028 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_31_603
timestamp 1644511149
transform 1 0 56580 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_31_615
timestamp 1644511149
transform 1 0 57684 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_620
timestamp 1644511149
transform 1 0 58144 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_624
timestamp 1644511149
transform 1 0 58512 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_3
timestamp 1644511149
transform 1 0 1380 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_15
timestamp 1644511149
transform 1 0 2484 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_27
timestamp 1644511149
transform 1 0 3588 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_29
timestamp 1644511149
transform 1 0 3772 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_41
timestamp 1644511149
transform 1 0 4876 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_53
timestamp 1644511149
transform 1 0 5980 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_65
timestamp 1644511149
transform 1 0 7084 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_77
timestamp 1644511149
transform 1 0 8188 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_83
timestamp 1644511149
transform 1 0 8740 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_85
timestamp 1644511149
transform 1 0 8924 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_97
timestamp 1644511149
transform 1 0 10028 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_109
timestamp 1644511149
transform 1 0 11132 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_121
timestamp 1644511149
transform 1 0 12236 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_133
timestamp 1644511149
transform 1 0 13340 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_139
timestamp 1644511149
transform 1 0 13892 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_141
timestamp 1644511149
transform 1 0 14076 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_153
timestamp 1644511149
transform 1 0 15180 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_165
timestamp 1644511149
transform 1 0 16284 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_177
timestamp 1644511149
transform 1 0 17388 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_189
timestamp 1644511149
transform 1 0 18492 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_195
timestamp 1644511149
transform 1 0 19044 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_197
timestamp 1644511149
transform 1 0 19228 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_209
timestamp 1644511149
transform 1 0 20332 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_221
timestamp 1644511149
transform 1 0 21436 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_233
timestamp 1644511149
transform 1 0 22540 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_245
timestamp 1644511149
transform 1 0 23644 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_251
timestamp 1644511149
transform 1 0 24196 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_253
timestamp 1644511149
transform 1 0 24380 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_265
timestamp 1644511149
transform 1 0 25484 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_277
timestamp 1644511149
transform 1 0 26588 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_289
timestamp 1644511149
transform 1 0 27692 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_301
timestamp 1644511149
transform 1 0 28796 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_307
timestamp 1644511149
transform 1 0 29348 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_309
timestamp 1644511149
transform 1 0 29532 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_321
timestamp 1644511149
transform 1 0 30636 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_333
timestamp 1644511149
transform 1 0 31740 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_345
timestamp 1644511149
transform 1 0 32844 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_357
timestamp 1644511149
transform 1 0 33948 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_363
timestamp 1644511149
transform 1 0 34500 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_365
timestamp 1644511149
transform 1 0 34684 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_377
timestamp 1644511149
transform 1 0 35788 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_389
timestamp 1644511149
transform 1 0 36892 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_401
timestamp 1644511149
transform 1 0 37996 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_413
timestamp 1644511149
transform 1 0 39100 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_419
timestamp 1644511149
transform 1 0 39652 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_421
timestamp 1644511149
transform 1 0 39836 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_433
timestamp 1644511149
transform 1 0 40940 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_445
timestamp 1644511149
transform 1 0 42044 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_457
timestamp 1644511149
transform 1 0 43148 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_469
timestamp 1644511149
transform 1 0 44252 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_475
timestamp 1644511149
transform 1 0 44804 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_477
timestamp 1644511149
transform 1 0 44988 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_489
timestamp 1644511149
transform 1 0 46092 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_501
timestamp 1644511149
transform 1 0 47196 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_513
timestamp 1644511149
transform 1 0 48300 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_525
timestamp 1644511149
transform 1 0 49404 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_531
timestamp 1644511149
transform 1 0 49956 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_533
timestamp 1644511149
transform 1 0 50140 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_545
timestamp 1644511149
transform 1 0 51244 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_557
timestamp 1644511149
transform 1 0 52348 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_569
timestamp 1644511149
transform 1 0 53452 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_581
timestamp 1644511149
transform 1 0 54556 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_587
timestamp 1644511149
transform 1 0 55108 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_589
timestamp 1644511149
transform 1 0 55292 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_601
timestamp 1644511149
transform 1 0 56396 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_613
timestamp 1644511149
transform 1 0 57500 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_3
timestamp 1644511149
transform 1 0 1380 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_15
timestamp 1644511149
transform 1 0 2484 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_27
timestamp 1644511149
transform 1 0 3588 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_39
timestamp 1644511149
transform 1 0 4692 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_51
timestamp 1644511149
transform 1 0 5796 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_55
timestamp 1644511149
transform 1 0 6164 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_57
timestamp 1644511149
transform 1 0 6348 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_69
timestamp 1644511149
transform 1 0 7452 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_81
timestamp 1644511149
transform 1 0 8556 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_93
timestamp 1644511149
transform 1 0 9660 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_105
timestamp 1644511149
transform 1 0 10764 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_111
timestamp 1644511149
transform 1 0 11316 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_113
timestamp 1644511149
transform 1 0 11500 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_125
timestamp 1644511149
transform 1 0 12604 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_137
timestamp 1644511149
transform 1 0 13708 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_149
timestamp 1644511149
transform 1 0 14812 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_161
timestamp 1644511149
transform 1 0 15916 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_167
timestamp 1644511149
transform 1 0 16468 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_169
timestamp 1644511149
transform 1 0 16652 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_181
timestamp 1644511149
transform 1 0 17756 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_193
timestamp 1644511149
transform 1 0 18860 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_205
timestamp 1644511149
transform 1 0 19964 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_217
timestamp 1644511149
transform 1 0 21068 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_223
timestamp 1644511149
transform 1 0 21620 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_225
timestamp 1644511149
transform 1 0 21804 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_237
timestamp 1644511149
transform 1 0 22908 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_249
timestamp 1644511149
transform 1 0 24012 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_261
timestamp 1644511149
transform 1 0 25116 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_273
timestamp 1644511149
transform 1 0 26220 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_279
timestamp 1644511149
transform 1 0 26772 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_281
timestamp 1644511149
transform 1 0 26956 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_293
timestamp 1644511149
transform 1 0 28060 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_305
timestamp 1644511149
transform 1 0 29164 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_317
timestamp 1644511149
transform 1 0 30268 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_329
timestamp 1644511149
transform 1 0 31372 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_335
timestamp 1644511149
transform 1 0 31924 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_337
timestamp 1644511149
transform 1 0 32108 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_349
timestamp 1644511149
transform 1 0 33212 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_361
timestamp 1644511149
transform 1 0 34316 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_373
timestamp 1644511149
transform 1 0 35420 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_385
timestamp 1644511149
transform 1 0 36524 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_391
timestamp 1644511149
transform 1 0 37076 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_393
timestamp 1644511149
transform 1 0 37260 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_405
timestamp 1644511149
transform 1 0 38364 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_417
timestamp 1644511149
transform 1 0 39468 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_429
timestamp 1644511149
transform 1 0 40572 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_441
timestamp 1644511149
transform 1 0 41676 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_447
timestamp 1644511149
transform 1 0 42228 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_449
timestamp 1644511149
transform 1 0 42412 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_461
timestamp 1644511149
transform 1 0 43516 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_473
timestamp 1644511149
transform 1 0 44620 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_485
timestamp 1644511149
transform 1 0 45724 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_497
timestamp 1644511149
transform 1 0 46828 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_503
timestamp 1644511149
transform 1 0 47380 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_505
timestamp 1644511149
transform 1 0 47564 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_517
timestamp 1644511149
transform 1 0 48668 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_529
timestamp 1644511149
transform 1 0 49772 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_541
timestamp 1644511149
transform 1 0 50876 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_553
timestamp 1644511149
transform 1 0 51980 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_559
timestamp 1644511149
transform 1 0 52532 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_561
timestamp 1644511149
transform 1 0 52716 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_573
timestamp 1644511149
transform 1 0 53820 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_585
timestamp 1644511149
transform 1 0 54924 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_597
timestamp 1644511149
transform 1 0 56028 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_609
timestamp 1644511149
transform 1 0 57132 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_615
timestamp 1644511149
transform 1 0 57684 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_617
timestamp 1644511149
transform 1 0 57868 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_34_3
timestamp 1644511149
transform 1 0 1380 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_15
timestamp 1644511149
transform 1 0 2484 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_27
timestamp 1644511149
transform 1 0 3588 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_29
timestamp 1644511149
transform 1 0 3772 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_41
timestamp 1644511149
transform 1 0 4876 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_53
timestamp 1644511149
transform 1 0 5980 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_65
timestamp 1644511149
transform 1 0 7084 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_77
timestamp 1644511149
transform 1 0 8188 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_83
timestamp 1644511149
transform 1 0 8740 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_85
timestamp 1644511149
transform 1 0 8924 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_97
timestamp 1644511149
transform 1 0 10028 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_109
timestamp 1644511149
transform 1 0 11132 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_121
timestamp 1644511149
transform 1 0 12236 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_133
timestamp 1644511149
transform 1 0 13340 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_139
timestamp 1644511149
transform 1 0 13892 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_141
timestamp 1644511149
transform 1 0 14076 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_153
timestamp 1644511149
transform 1 0 15180 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_165
timestamp 1644511149
transform 1 0 16284 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_177
timestamp 1644511149
transform 1 0 17388 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_189
timestamp 1644511149
transform 1 0 18492 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_195
timestamp 1644511149
transform 1 0 19044 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_197
timestamp 1644511149
transform 1 0 19228 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_209
timestamp 1644511149
transform 1 0 20332 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_221
timestamp 1644511149
transform 1 0 21436 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_233
timestamp 1644511149
transform 1 0 22540 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_245
timestamp 1644511149
transform 1 0 23644 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_251
timestamp 1644511149
transform 1 0 24196 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_253
timestamp 1644511149
transform 1 0 24380 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_265
timestamp 1644511149
transform 1 0 25484 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_277
timestamp 1644511149
transform 1 0 26588 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_289
timestamp 1644511149
transform 1 0 27692 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_301
timestamp 1644511149
transform 1 0 28796 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_307
timestamp 1644511149
transform 1 0 29348 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_309
timestamp 1644511149
transform 1 0 29532 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_321
timestamp 1644511149
transform 1 0 30636 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_333
timestamp 1644511149
transform 1 0 31740 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_345
timestamp 1644511149
transform 1 0 32844 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_357
timestamp 1644511149
transform 1 0 33948 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_363
timestamp 1644511149
transform 1 0 34500 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_365
timestamp 1644511149
transform 1 0 34684 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_377
timestamp 1644511149
transform 1 0 35788 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_389
timestamp 1644511149
transform 1 0 36892 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_401
timestamp 1644511149
transform 1 0 37996 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_413
timestamp 1644511149
transform 1 0 39100 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_419
timestamp 1644511149
transform 1 0 39652 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_421
timestamp 1644511149
transform 1 0 39836 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_433
timestamp 1644511149
transform 1 0 40940 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_445
timestamp 1644511149
transform 1 0 42044 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_457
timestamp 1644511149
transform 1 0 43148 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_469
timestamp 1644511149
transform 1 0 44252 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_475
timestamp 1644511149
transform 1 0 44804 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_477
timestamp 1644511149
transform 1 0 44988 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_489
timestamp 1644511149
transform 1 0 46092 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_501
timestamp 1644511149
transform 1 0 47196 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_513
timestamp 1644511149
transform 1 0 48300 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_525
timestamp 1644511149
transform 1 0 49404 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_531
timestamp 1644511149
transform 1 0 49956 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_533
timestamp 1644511149
transform 1 0 50140 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_545
timestamp 1644511149
transform 1 0 51244 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_557
timestamp 1644511149
transform 1 0 52348 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_569
timestamp 1644511149
transform 1 0 53452 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_581
timestamp 1644511149
transform 1 0 54556 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_587
timestamp 1644511149
transform 1 0 55108 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_589
timestamp 1644511149
transform 1 0 55292 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_601
timestamp 1644511149
transform 1 0 56396 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_613
timestamp 1644511149
transform 1 0 57500 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_3
timestamp 1644511149
transform 1 0 1380 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_15
timestamp 1644511149
transform 1 0 2484 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_27
timestamp 1644511149
transform 1 0 3588 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_39
timestamp 1644511149
transform 1 0 4692 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_51
timestamp 1644511149
transform 1 0 5796 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_55
timestamp 1644511149
transform 1 0 6164 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_57
timestamp 1644511149
transform 1 0 6348 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_69
timestamp 1644511149
transform 1 0 7452 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_81
timestamp 1644511149
transform 1 0 8556 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_93
timestamp 1644511149
transform 1 0 9660 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_105
timestamp 1644511149
transform 1 0 10764 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_111
timestamp 1644511149
transform 1 0 11316 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_113
timestamp 1644511149
transform 1 0 11500 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_125
timestamp 1644511149
transform 1 0 12604 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_137
timestamp 1644511149
transform 1 0 13708 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_149
timestamp 1644511149
transform 1 0 14812 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_161
timestamp 1644511149
transform 1 0 15916 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_167
timestamp 1644511149
transform 1 0 16468 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_169
timestamp 1644511149
transform 1 0 16652 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_181
timestamp 1644511149
transform 1 0 17756 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_193
timestamp 1644511149
transform 1 0 18860 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_205
timestamp 1644511149
transform 1 0 19964 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_217
timestamp 1644511149
transform 1 0 21068 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_223
timestamp 1644511149
transform 1 0 21620 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_225
timestamp 1644511149
transform 1 0 21804 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_237
timestamp 1644511149
transform 1 0 22908 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_249
timestamp 1644511149
transform 1 0 24012 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_261
timestamp 1644511149
transform 1 0 25116 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_273
timestamp 1644511149
transform 1 0 26220 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_279
timestamp 1644511149
transform 1 0 26772 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_281
timestamp 1644511149
transform 1 0 26956 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_293
timestamp 1644511149
transform 1 0 28060 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_305
timestamp 1644511149
transform 1 0 29164 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_317
timestamp 1644511149
transform 1 0 30268 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_329
timestamp 1644511149
transform 1 0 31372 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_335
timestamp 1644511149
transform 1 0 31924 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_337
timestamp 1644511149
transform 1 0 32108 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_349
timestamp 1644511149
transform 1 0 33212 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_361
timestamp 1644511149
transform 1 0 34316 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_373
timestamp 1644511149
transform 1 0 35420 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_385
timestamp 1644511149
transform 1 0 36524 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_391
timestamp 1644511149
transform 1 0 37076 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_393
timestamp 1644511149
transform 1 0 37260 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_405
timestamp 1644511149
transform 1 0 38364 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_417
timestamp 1644511149
transform 1 0 39468 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_429
timestamp 1644511149
transform 1 0 40572 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_441
timestamp 1644511149
transform 1 0 41676 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_447
timestamp 1644511149
transform 1 0 42228 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_449
timestamp 1644511149
transform 1 0 42412 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_461
timestamp 1644511149
transform 1 0 43516 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_473
timestamp 1644511149
transform 1 0 44620 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_485
timestamp 1644511149
transform 1 0 45724 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_497
timestamp 1644511149
transform 1 0 46828 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_503
timestamp 1644511149
transform 1 0 47380 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_505
timestamp 1644511149
transform 1 0 47564 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_517
timestamp 1644511149
transform 1 0 48668 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_529
timestamp 1644511149
transform 1 0 49772 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_541
timestamp 1644511149
transform 1 0 50876 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_553
timestamp 1644511149
transform 1 0 51980 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_559
timestamp 1644511149
transform 1 0 52532 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_561
timestamp 1644511149
transform 1 0 52716 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_573
timestamp 1644511149
transform 1 0 53820 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_585
timestamp 1644511149
transform 1 0 54924 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_597
timestamp 1644511149
transform 1 0 56028 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_609
timestamp 1644511149
transform 1 0 57132 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_615
timestamp 1644511149
transform 1 0 57684 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_35_617
timestamp 1644511149
transform 1 0 57868 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_36_3
timestamp 1644511149
transform 1 0 1380 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_15
timestamp 1644511149
transform 1 0 2484 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_27
timestamp 1644511149
transform 1 0 3588 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_29
timestamp 1644511149
transform 1 0 3772 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_41
timestamp 1644511149
transform 1 0 4876 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_53
timestamp 1644511149
transform 1 0 5980 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_65
timestamp 1644511149
transform 1 0 7084 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_77
timestamp 1644511149
transform 1 0 8188 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_83
timestamp 1644511149
transform 1 0 8740 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_85
timestamp 1644511149
transform 1 0 8924 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_97
timestamp 1644511149
transform 1 0 10028 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_109
timestamp 1644511149
transform 1 0 11132 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_121
timestamp 1644511149
transform 1 0 12236 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_133
timestamp 1644511149
transform 1 0 13340 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_139
timestamp 1644511149
transform 1 0 13892 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_141
timestamp 1644511149
transform 1 0 14076 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_153
timestamp 1644511149
transform 1 0 15180 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_165
timestamp 1644511149
transform 1 0 16284 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_177
timestamp 1644511149
transform 1 0 17388 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_189
timestamp 1644511149
transform 1 0 18492 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_195
timestamp 1644511149
transform 1 0 19044 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_197
timestamp 1644511149
transform 1 0 19228 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_209
timestamp 1644511149
transform 1 0 20332 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_221
timestamp 1644511149
transform 1 0 21436 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_233
timestamp 1644511149
transform 1 0 22540 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_245
timestamp 1644511149
transform 1 0 23644 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_251
timestamp 1644511149
transform 1 0 24196 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_253
timestamp 1644511149
transform 1 0 24380 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_265
timestamp 1644511149
transform 1 0 25484 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_277
timestamp 1644511149
transform 1 0 26588 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_289
timestamp 1644511149
transform 1 0 27692 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_301
timestamp 1644511149
transform 1 0 28796 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_307
timestamp 1644511149
transform 1 0 29348 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_309
timestamp 1644511149
transform 1 0 29532 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_321
timestamp 1644511149
transform 1 0 30636 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_333
timestamp 1644511149
transform 1 0 31740 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_345
timestamp 1644511149
transform 1 0 32844 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_357
timestamp 1644511149
transform 1 0 33948 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_363
timestamp 1644511149
transform 1 0 34500 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_365
timestamp 1644511149
transform 1 0 34684 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_377
timestamp 1644511149
transform 1 0 35788 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_389
timestamp 1644511149
transform 1 0 36892 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_401
timestamp 1644511149
transform 1 0 37996 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_413
timestamp 1644511149
transform 1 0 39100 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_419
timestamp 1644511149
transform 1 0 39652 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_421
timestamp 1644511149
transform 1 0 39836 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_433
timestamp 1644511149
transform 1 0 40940 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_445
timestamp 1644511149
transform 1 0 42044 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_457
timestamp 1644511149
transform 1 0 43148 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_469
timestamp 1644511149
transform 1 0 44252 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_475
timestamp 1644511149
transform 1 0 44804 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_477
timestamp 1644511149
transform 1 0 44988 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_489
timestamp 1644511149
transform 1 0 46092 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_501
timestamp 1644511149
transform 1 0 47196 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_513
timestamp 1644511149
transform 1 0 48300 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_525
timestamp 1644511149
transform 1 0 49404 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_531
timestamp 1644511149
transform 1 0 49956 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_533
timestamp 1644511149
transform 1 0 50140 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_545
timestamp 1644511149
transform 1 0 51244 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_557
timestamp 1644511149
transform 1 0 52348 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_569
timestamp 1644511149
transform 1 0 53452 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_581
timestamp 1644511149
transform 1 0 54556 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_587
timestamp 1644511149
transform 1 0 55108 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_589
timestamp 1644511149
transform 1 0 55292 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_601
timestamp 1644511149
transform 1 0 56396 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_613
timestamp 1644511149
transform 1 0 57500 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_3
timestamp 1644511149
transform 1 0 1380 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_15
timestamp 1644511149
transform 1 0 2484 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_27
timestamp 1644511149
transform 1 0 3588 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_39
timestamp 1644511149
transform 1 0 4692 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_51
timestamp 1644511149
transform 1 0 5796 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_55
timestamp 1644511149
transform 1 0 6164 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_57
timestamp 1644511149
transform 1 0 6348 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_37_69
timestamp 1644511149
transform 1 0 7452 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_90
timestamp 1644511149
transform 1 0 9384 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_102
timestamp 1644511149
transform 1 0 10488 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_37_110
timestamp 1644511149
transform 1 0 11224 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_37_113
timestamp 1644511149
transform 1 0 11500 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_125
timestamp 1644511149
transform 1 0 12604 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_137
timestamp 1644511149
transform 1 0 13708 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_149
timestamp 1644511149
transform 1 0 14812 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_161
timestamp 1644511149
transform 1 0 15916 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_167
timestamp 1644511149
transform 1 0 16468 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_169
timestamp 1644511149
transform 1 0 16652 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_181
timestamp 1644511149
transform 1 0 17756 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_193
timestamp 1644511149
transform 1 0 18860 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_205
timestamp 1644511149
transform 1 0 19964 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_217
timestamp 1644511149
transform 1 0 21068 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_223
timestamp 1644511149
transform 1 0 21620 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_225
timestamp 1644511149
transform 1 0 21804 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_237
timestamp 1644511149
transform 1 0 22908 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_249
timestamp 1644511149
transform 1 0 24012 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_261
timestamp 1644511149
transform 1 0 25116 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_273
timestamp 1644511149
transform 1 0 26220 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_279
timestamp 1644511149
transform 1 0 26772 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_281
timestamp 1644511149
transform 1 0 26956 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_293
timestamp 1644511149
transform 1 0 28060 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_305
timestamp 1644511149
transform 1 0 29164 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_317
timestamp 1644511149
transform 1 0 30268 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_329
timestamp 1644511149
transform 1 0 31372 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_335
timestamp 1644511149
transform 1 0 31924 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_337
timestamp 1644511149
transform 1 0 32108 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_349
timestamp 1644511149
transform 1 0 33212 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_361
timestamp 1644511149
transform 1 0 34316 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_373
timestamp 1644511149
transform 1 0 35420 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_385
timestamp 1644511149
transform 1 0 36524 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_391
timestamp 1644511149
transform 1 0 37076 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_393
timestamp 1644511149
transform 1 0 37260 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_405
timestamp 1644511149
transform 1 0 38364 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_417
timestamp 1644511149
transform 1 0 39468 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_429
timestamp 1644511149
transform 1 0 40572 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_441
timestamp 1644511149
transform 1 0 41676 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_447
timestamp 1644511149
transform 1 0 42228 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_449
timestamp 1644511149
transform 1 0 42412 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_461
timestamp 1644511149
transform 1 0 43516 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_473
timestamp 1644511149
transform 1 0 44620 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_485
timestamp 1644511149
transform 1 0 45724 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_497
timestamp 1644511149
transform 1 0 46828 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_503
timestamp 1644511149
transform 1 0 47380 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_505
timestamp 1644511149
transform 1 0 47564 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_517
timestamp 1644511149
transform 1 0 48668 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_529
timestamp 1644511149
transform 1 0 49772 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_541
timestamp 1644511149
transform 1 0 50876 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_553
timestamp 1644511149
transform 1 0 51980 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_559
timestamp 1644511149
transform 1 0 52532 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_561
timestamp 1644511149
transform 1 0 52716 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_573
timestamp 1644511149
transform 1 0 53820 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_585
timestamp 1644511149
transform 1 0 54924 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_597
timestamp 1644511149
transform 1 0 56028 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_609
timestamp 1644511149
transform 1 0 57132 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_615
timestamp 1644511149
transform 1 0 57684 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_37_617
timestamp 1644511149
transform 1 0 57868 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_38_3
timestamp 1644511149
transform 1 0 1380 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_15
timestamp 1644511149
transform 1 0 2484 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_38_27
timestamp 1644511149
transform 1 0 3588 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_29
timestamp 1644511149
transform 1 0 3772 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_41
timestamp 1644511149
transform 1 0 4876 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_53
timestamp 1644511149
transform 1 0 5980 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_65
timestamp 1644511149
transform 1 0 7084 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_38_80
timestamp 1644511149
transform 1 0 8464 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_38_85
timestamp 1644511149
transform 1 0 8924 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_97
timestamp 1644511149
transform 1 0 10028 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_109
timestamp 1644511149
transform 1 0 11132 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_121
timestamp 1644511149
transform 1 0 12236 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_133
timestamp 1644511149
transform 1 0 13340 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_139
timestamp 1644511149
transform 1 0 13892 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_141
timestamp 1644511149
transform 1 0 14076 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_153
timestamp 1644511149
transform 1 0 15180 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_165
timestamp 1644511149
transform 1 0 16284 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_177
timestamp 1644511149
transform 1 0 17388 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_189
timestamp 1644511149
transform 1 0 18492 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_195
timestamp 1644511149
transform 1 0 19044 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_197
timestamp 1644511149
transform 1 0 19228 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_209
timestamp 1644511149
transform 1 0 20332 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_221
timestamp 1644511149
transform 1 0 21436 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_233
timestamp 1644511149
transform 1 0 22540 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_245
timestamp 1644511149
transform 1 0 23644 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_251
timestamp 1644511149
transform 1 0 24196 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_253
timestamp 1644511149
transform 1 0 24380 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_265
timestamp 1644511149
transform 1 0 25484 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_277
timestamp 1644511149
transform 1 0 26588 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_289
timestamp 1644511149
transform 1 0 27692 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_301
timestamp 1644511149
transform 1 0 28796 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_307
timestamp 1644511149
transform 1 0 29348 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_309
timestamp 1644511149
transform 1 0 29532 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_321
timestamp 1644511149
transform 1 0 30636 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_333
timestamp 1644511149
transform 1 0 31740 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_345
timestamp 1644511149
transform 1 0 32844 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_357
timestamp 1644511149
transform 1 0 33948 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_363
timestamp 1644511149
transform 1 0 34500 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_365
timestamp 1644511149
transform 1 0 34684 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_377
timestamp 1644511149
transform 1 0 35788 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_389
timestamp 1644511149
transform 1 0 36892 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_401
timestamp 1644511149
transform 1 0 37996 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_413
timestamp 1644511149
transform 1 0 39100 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_419
timestamp 1644511149
transform 1 0 39652 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_421
timestamp 1644511149
transform 1 0 39836 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_433
timestamp 1644511149
transform 1 0 40940 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_445
timestamp 1644511149
transform 1 0 42044 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_457
timestamp 1644511149
transform 1 0 43148 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_469
timestamp 1644511149
transform 1 0 44252 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_475
timestamp 1644511149
transform 1 0 44804 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_477
timestamp 1644511149
transform 1 0 44988 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_489
timestamp 1644511149
transform 1 0 46092 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_501
timestamp 1644511149
transform 1 0 47196 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_513
timestamp 1644511149
transform 1 0 48300 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_525
timestamp 1644511149
transform 1 0 49404 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_531
timestamp 1644511149
transform 1 0 49956 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_533
timestamp 1644511149
transform 1 0 50140 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_545
timestamp 1644511149
transform 1 0 51244 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_557
timestamp 1644511149
transform 1 0 52348 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_569
timestamp 1644511149
transform 1 0 53452 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_581
timestamp 1644511149
transform 1 0 54556 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_587
timestamp 1644511149
transform 1 0 55108 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_589
timestamp 1644511149
transform 1 0 55292 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_601
timestamp 1644511149
transform 1 0 56396 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_613
timestamp 1644511149
transform 1 0 57500 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_3
timestamp 1644511149
transform 1 0 1380 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_15
timestamp 1644511149
transform 1 0 2484 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_27
timestamp 1644511149
transform 1 0 3588 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_39
timestamp 1644511149
transform 1 0 4692 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_51
timestamp 1644511149
transform 1 0 5796 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_55
timestamp 1644511149
transform 1 0 6164 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_57
timestamp 1644511149
transform 1 0 6348 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_69
timestamp 1644511149
transform 1 0 7452 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_81
timestamp 1644511149
transform 1 0 8556 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_93
timestamp 1644511149
transform 1 0 9660 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_105
timestamp 1644511149
transform 1 0 10764 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_111
timestamp 1644511149
transform 1 0 11316 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_113
timestamp 1644511149
transform 1 0 11500 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_125
timestamp 1644511149
transform 1 0 12604 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_137
timestamp 1644511149
transform 1 0 13708 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_149
timestamp 1644511149
transform 1 0 14812 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_161
timestamp 1644511149
transform 1 0 15916 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_167
timestamp 1644511149
transform 1 0 16468 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_169
timestamp 1644511149
transform 1 0 16652 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_181
timestamp 1644511149
transform 1 0 17756 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_193
timestamp 1644511149
transform 1 0 18860 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_205
timestamp 1644511149
transform 1 0 19964 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_217
timestamp 1644511149
transform 1 0 21068 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_223
timestamp 1644511149
transform 1 0 21620 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_225
timestamp 1644511149
transform 1 0 21804 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_237
timestamp 1644511149
transform 1 0 22908 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_249
timestamp 1644511149
transform 1 0 24012 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_261
timestamp 1644511149
transform 1 0 25116 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_273
timestamp 1644511149
transform 1 0 26220 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_279
timestamp 1644511149
transform 1 0 26772 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_281
timestamp 1644511149
transform 1 0 26956 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_293
timestamp 1644511149
transform 1 0 28060 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_305
timestamp 1644511149
transform 1 0 29164 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_317
timestamp 1644511149
transform 1 0 30268 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_329
timestamp 1644511149
transform 1 0 31372 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_335
timestamp 1644511149
transform 1 0 31924 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_337
timestamp 1644511149
transform 1 0 32108 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_349
timestamp 1644511149
transform 1 0 33212 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_361
timestamp 1644511149
transform 1 0 34316 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_373
timestamp 1644511149
transform 1 0 35420 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_385
timestamp 1644511149
transform 1 0 36524 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_391
timestamp 1644511149
transform 1 0 37076 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_393
timestamp 1644511149
transform 1 0 37260 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_405
timestamp 1644511149
transform 1 0 38364 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_417
timestamp 1644511149
transform 1 0 39468 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_429
timestamp 1644511149
transform 1 0 40572 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_441
timestamp 1644511149
transform 1 0 41676 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_447
timestamp 1644511149
transform 1 0 42228 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_449
timestamp 1644511149
transform 1 0 42412 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_461
timestamp 1644511149
transform 1 0 43516 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_473
timestamp 1644511149
transform 1 0 44620 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_485
timestamp 1644511149
transform 1 0 45724 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_497
timestamp 1644511149
transform 1 0 46828 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_503
timestamp 1644511149
transform 1 0 47380 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_505
timestamp 1644511149
transform 1 0 47564 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_517
timestamp 1644511149
transform 1 0 48668 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_529
timestamp 1644511149
transform 1 0 49772 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_541
timestamp 1644511149
transform 1 0 50876 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_553
timestamp 1644511149
transform 1 0 51980 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_559
timestamp 1644511149
transform 1 0 52532 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_561
timestamp 1644511149
transform 1 0 52716 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_573
timestamp 1644511149
transform 1 0 53820 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_585
timestamp 1644511149
transform 1 0 54924 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_39_609
timestamp 1644511149
transform 1 0 57132 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_615
timestamp 1644511149
transform 1 0 57684 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_39_617
timestamp 1644511149
transform 1 0 57868 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_40_3
timestamp 1644511149
transform 1 0 1380 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_15
timestamp 1644511149
transform 1 0 2484 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_27
timestamp 1644511149
transform 1 0 3588 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_29
timestamp 1644511149
transform 1 0 3772 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_41
timestamp 1644511149
transform 1 0 4876 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_53
timestamp 1644511149
transform 1 0 5980 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_65
timestamp 1644511149
transform 1 0 7084 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_77
timestamp 1644511149
transform 1 0 8188 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_83
timestamp 1644511149
transform 1 0 8740 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_85
timestamp 1644511149
transform 1 0 8924 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_97
timestamp 1644511149
transform 1 0 10028 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_109
timestamp 1644511149
transform 1 0 11132 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_121
timestamp 1644511149
transform 1 0 12236 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_133
timestamp 1644511149
transform 1 0 13340 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_139
timestamp 1644511149
transform 1 0 13892 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_141
timestamp 1644511149
transform 1 0 14076 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_153
timestamp 1644511149
transform 1 0 15180 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_165
timestamp 1644511149
transform 1 0 16284 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_177
timestamp 1644511149
transform 1 0 17388 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_189
timestamp 1644511149
transform 1 0 18492 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_195
timestamp 1644511149
transform 1 0 19044 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_197
timestamp 1644511149
transform 1 0 19228 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_209
timestamp 1644511149
transform 1 0 20332 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_221
timestamp 1644511149
transform 1 0 21436 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_233
timestamp 1644511149
transform 1 0 22540 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_245
timestamp 1644511149
transform 1 0 23644 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_251
timestamp 1644511149
transform 1 0 24196 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_253
timestamp 1644511149
transform 1 0 24380 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_265
timestamp 1644511149
transform 1 0 25484 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_277
timestamp 1644511149
transform 1 0 26588 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_289
timestamp 1644511149
transform 1 0 27692 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_301
timestamp 1644511149
transform 1 0 28796 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_307
timestamp 1644511149
transform 1 0 29348 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_309
timestamp 1644511149
transform 1 0 29532 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_321
timestamp 1644511149
transform 1 0 30636 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_333
timestamp 1644511149
transform 1 0 31740 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_345
timestamp 1644511149
transform 1 0 32844 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_357
timestamp 1644511149
transform 1 0 33948 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_363
timestamp 1644511149
transform 1 0 34500 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_365
timestamp 1644511149
transform 1 0 34684 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_377
timestamp 1644511149
transform 1 0 35788 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_389
timestamp 1644511149
transform 1 0 36892 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_401
timestamp 1644511149
transform 1 0 37996 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_413
timestamp 1644511149
transform 1 0 39100 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_419
timestamp 1644511149
transform 1 0 39652 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_421
timestamp 1644511149
transform 1 0 39836 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_433
timestamp 1644511149
transform 1 0 40940 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_445
timestamp 1644511149
transform 1 0 42044 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_457
timestamp 1644511149
transform 1 0 43148 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_469
timestamp 1644511149
transform 1 0 44252 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_475
timestamp 1644511149
transform 1 0 44804 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_477
timestamp 1644511149
transform 1 0 44988 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_489
timestamp 1644511149
transform 1 0 46092 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_501
timestamp 1644511149
transform 1 0 47196 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_513
timestamp 1644511149
transform 1 0 48300 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_525
timestamp 1644511149
transform 1 0 49404 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_531
timestamp 1644511149
transform 1 0 49956 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_533
timestamp 1644511149
transform 1 0 50140 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_545
timestamp 1644511149
transform 1 0 51244 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_557
timestamp 1644511149
transform 1 0 52348 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_569
timestamp 1644511149
transform 1 0 53452 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_581
timestamp 1644511149
transform 1 0 54556 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_587
timestamp 1644511149
transform 1 0 55108 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_40_589
timestamp 1644511149
transform 1 0 55292 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_40_597
timestamp 1644511149
transform 1 0 56028 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_40_621
timestamp 1644511149
transform 1 0 58236 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_41_3
timestamp 1644511149
transform 1 0 1380 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_15
timestamp 1644511149
transform 1 0 2484 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_27
timestamp 1644511149
transform 1 0 3588 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_39
timestamp 1644511149
transform 1 0 4692 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_51
timestamp 1644511149
transform 1 0 5796 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_55
timestamp 1644511149
transform 1 0 6164 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_57
timestamp 1644511149
transform 1 0 6348 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_69
timestamp 1644511149
transform 1 0 7452 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_41_81
timestamp 1644511149
transform 1 0 8556 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_41_99
timestamp 1644511149
transform 1 0 10212 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_41_111
timestamp 1644511149
transform 1 0 11316 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_113
timestamp 1644511149
transform 1 0 11500 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_125
timestamp 1644511149
transform 1 0 12604 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_137
timestamp 1644511149
transform 1 0 13708 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_149
timestamp 1644511149
transform 1 0 14812 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_161
timestamp 1644511149
transform 1 0 15916 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_167
timestamp 1644511149
transform 1 0 16468 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_169
timestamp 1644511149
transform 1 0 16652 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_181
timestamp 1644511149
transform 1 0 17756 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_193
timestamp 1644511149
transform 1 0 18860 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_205
timestamp 1644511149
transform 1 0 19964 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_217
timestamp 1644511149
transform 1 0 21068 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_223
timestamp 1644511149
transform 1 0 21620 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_225
timestamp 1644511149
transform 1 0 21804 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_237
timestamp 1644511149
transform 1 0 22908 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_249
timestamp 1644511149
transform 1 0 24012 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_261
timestamp 1644511149
transform 1 0 25116 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_273
timestamp 1644511149
transform 1 0 26220 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_279
timestamp 1644511149
transform 1 0 26772 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_281
timestamp 1644511149
transform 1 0 26956 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_293
timestamp 1644511149
transform 1 0 28060 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_305
timestamp 1644511149
transform 1 0 29164 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_317
timestamp 1644511149
transform 1 0 30268 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_329
timestamp 1644511149
transform 1 0 31372 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_335
timestamp 1644511149
transform 1 0 31924 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_337
timestamp 1644511149
transform 1 0 32108 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_349
timestamp 1644511149
transform 1 0 33212 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_361
timestamp 1644511149
transform 1 0 34316 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_373
timestamp 1644511149
transform 1 0 35420 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_385
timestamp 1644511149
transform 1 0 36524 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_391
timestamp 1644511149
transform 1 0 37076 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_393
timestamp 1644511149
transform 1 0 37260 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_405
timestamp 1644511149
transform 1 0 38364 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_417
timestamp 1644511149
transform 1 0 39468 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_429
timestamp 1644511149
transform 1 0 40572 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_441
timestamp 1644511149
transform 1 0 41676 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_447
timestamp 1644511149
transform 1 0 42228 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_449
timestamp 1644511149
transform 1 0 42412 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_461
timestamp 1644511149
transform 1 0 43516 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_473
timestamp 1644511149
transform 1 0 44620 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_485
timestamp 1644511149
transform 1 0 45724 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_497
timestamp 1644511149
transform 1 0 46828 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_503
timestamp 1644511149
transform 1 0 47380 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_505
timestamp 1644511149
transform 1 0 47564 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_517
timestamp 1644511149
transform 1 0 48668 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_529
timestamp 1644511149
transform 1 0 49772 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_541
timestamp 1644511149
transform 1 0 50876 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_553
timestamp 1644511149
transform 1 0 51980 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_559
timestamp 1644511149
transform 1 0 52532 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_561
timestamp 1644511149
transform 1 0 52716 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_573
timestamp 1644511149
transform 1 0 53820 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_585
timestamp 1644511149
transform 1 0 54924 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_589
timestamp 1644511149
transform 1 0 55292 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_602
timestamp 1644511149
transform 1 0 56488 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_41_609
timestamp 1644511149
transform 1 0 57132 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_615
timestamp 1644511149
transform 1 0 57684 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_620
timestamp 1644511149
transform 1 0 58144 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_624
timestamp 1644511149
transform 1 0 58512 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_3
timestamp 1644511149
transform 1 0 1380 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_15
timestamp 1644511149
transform 1 0 2484 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_42_27
timestamp 1644511149
transform 1 0 3588 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_29
timestamp 1644511149
transform 1 0 3772 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_41
timestamp 1644511149
transform 1 0 4876 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_53
timestamp 1644511149
transform 1 0 5980 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_65
timestamp 1644511149
transform 1 0 7084 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_77
timestamp 1644511149
transform 1 0 8188 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_83
timestamp 1644511149
transform 1 0 8740 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_85
timestamp 1644511149
transform 1 0 8924 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_97
timestamp 1644511149
transform 1 0 10028 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_109
timestamp 1644511149
transform 1 0 11132 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_121
timestamp 1644511149
transform 1 0 12236 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_133
timestamp 1644511149
transform 1 0 13340 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_139
timestamp 1644511149
transform 1 0 13892 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_141
timestamp 1644511149
transform 1 0 14076 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_153
timestamp 1644511149
transform 1 0 15180 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_165
timestamp 1644511149
transform 1 0 16284 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_177
timestamp 1644511149
transform 1 0 17388 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_189
timestamp 1644511149
transform 1 0 18492 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_195
timestamp 1644511149
transform 1 0 19044 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_197
timestamp 1644511149
transform 1 0 19228 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_209
timestamp 1644511149
transform 1 0 20332 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_221
timestamp 1644511149
transform 1 0 21436 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_233
timestamp 1644511149
transform 1 0 22540 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_245
timestamp 1644511149
transform 1 0 23644 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_251
timestamp 1644511149
transform 1 0 24196 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_253
timestamp 1644511149
transform 1 0 24380 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_265
timestamp 1644511149
transform 1 0 25484 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_277
timestamp 1644511149
transform 1 0 26588 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_289
timestamp 1644511149
transform 1 0 27692 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_301
timestamp 1644511149
transform 1 0 28796 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_307
timestamp 1644511149
transform 1 0 29348 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_309
timestamp 1644511149
transform 1 0 29532 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_321
timestamp 1644511149
transform 1 0 30636 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_333
timestamp 1644511149
transform 1 0 31740 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_345
timestamp 1644511149
transform 1 0 32844 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_357
timestamp 1644511149
transform 1 0 33948 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_363
timestamp 1644511149
transform 1 0 34500 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_365
timestamp 1644511149
transform 1 0 34684 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_377
timestamp 1644511149
transform 1 0 35788 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_389
timestamp 1644511149
transform 1 0 36892 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_401
timestamp 1644511149
transform 1 0 37996 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_413
timestamp 1644511149
transform 1 0 39100 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_419
timestamp 1644511149
transform 1 0 39652 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_421
timestamp 1644511149
transform 1 0 39836 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_433
timestamp 1644511149
transform 1 0 40940 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_445
timestamp 1644511149
transform 1 0 42044 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_457
timestamp 1644511149
transform 1 0 43148 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_469
timestamp 1644511149
transform 1 0 44252 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_475
timestamp 1644511149
transform 1 0 44804 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_477
timestamp 1644511149
transform 1 0 44988 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_489
timestamp 1644511149
transform 1 0 46092 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_501
timestamp 1644511149
transform 1 0 47196 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_513
timestamp 1644511149
transform 1 0 48300 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_525
timestamp 1644511149
transform 1 0 49404 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_531
timestamp 1644511149
transform 1 0 49956 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_533
timestamp 1644511149
transform 1 0 50140 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_545
timestamp 1644511149
transform 1 0 51244 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_557
timestamp 1644511149
transform 1 0 52348 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_569
timestamp 1644511149
transform 1 0 53452 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_581
timestamp 1644511149
transform 1 0 54556 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_587
timestamp 1644511149
transform 1 0 55108 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_589
timestamp 1644511149
transform 1 0 55292 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_601
timestamp 1644511149
transform 1 0 56396 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_613
timestamp 1644511149
transform 1 0 57500 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_3
timestamp 1644511149
transform 1 0 1380 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_15
timestamp 1644511149
transform 1 0 2484 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_27
timestamp 1644511149
transform 1 0 3588 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_39
timestamp 1644511149
transform 1 0 4692 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_51
timestamp 1644511149
transform 1 0 5796 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_55
timestamp 1644511149
transform 1 0 6164 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_57
timestamp 1644511149
transform 1 0 6348 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_69
timestamp 1644511149
transform 1 0 7452 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_75
timestamp 1644511149
transform 1 0 8004 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_79
timestamp 1644511149
transform 1 0 8372 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_91
timestamp 1644511149
transform 1 0 9476 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_103
timestamp 1644511149
transform 1 0 10580 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_43_111
timestamp 1644511149
transform 1 0 11316 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_113
timestamp 1644511149
transform 1 0 11500 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_125
timestamp 1644511149
transform 1 0 12604 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_137
timestamp 1644511149
transform 1 0 13708 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_149
timestamp 1644511149
transform 1 0 14812 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_161
timestamp 1644511149
transform 1 0 15916 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_167
timestamp 1644511149
transform 1 0 16468 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_169
timestamp 1644511149
transform 1 0 16652 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_181
timestamp 1644511149
transform 1 0 17756 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_193
timestamp 1644511149
transform 1 0 18860 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_205
timestamp 1644511149
transform 1 0 19964 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_217
timestamp 1644511149
transform 1 0 21068 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_223
timestamp 1644511149
transform 1 0 21620 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_225
timestamp 1644511149
transform 1 0 21804 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_237
timestamp 1644511149
transform 1 0 22908 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_249
timestamp 1644511149
transform 1 0 24012 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_261
timestamp 1644511149
transform 1 0 25116 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_273
timestamp 1644511149
transform 1 0 26220 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_279
timestamp 1644511149
transform 1 0 26772 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_281
timestamp 1644511149
transform 1 0 26956 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_293
timestamp 1644511149
transform 1 0 28060 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_305
timestamp 1644511149
transform 1 0 29164 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_317
timestamp 1644511149
transform 1 0 30268 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_329
timestamp 1644511149
transform 1 0 31372 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_335
timestamp 1644511149
transform 1 0 31924 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_337
timestamp 1644511149
transform 1 0 32108 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_349
timestamp 1644511149
transform 1 0 33212 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_361
timestamp 1644511149
transform 1 0 34316 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_373
timestamp 1644511149
transform 1 0 35420 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_385
timestamp 1644511149
transform 1 0 36524 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_391
timestamp 1644511149
transform 1 0 37076 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_393
timestamp 1644511149
transform 1 0 37260 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_405
timestamp 1644511149
transform 1 0 38364 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_417
timestamp 1644511149
transform 1 0 39468 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_429
timestamp 1644511149
transform 1 0 40572 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_441
timestamp 1644511149
transform 1 0 41676 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_447
timestamp 1644511149
transform 1 0 42228 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_449
timestamp 1644511149
transform 1 0 42412 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_461
timestamp 1644511149
transform 1 0 43516 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_473
timestamp 1644511149
transform 1 0 44620 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_485
timestamp 1644511149
transform 1 0 45724 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_497
timestamp 1644511149
transform 1 0 46828 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_503
timestamp 1644511149
transform 1 0 47380 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_505
timestamp 1644511149
transform 1 0 47564 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_517
timestamp 1644511149
transform 1 0 48668 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_529
timestamp 1644511149
transform 1 0 49772 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_541
timestamp 1644511149
transform 1 0 50876 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_553
timestamp 1644511149
transform 1 0 51980 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_559
timestamp 1644511149
transform 1 0 52532 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_561
timestamp 1644511149
transform 1 0 52716 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_573
timestamp 1644511149
transform 1 0 53820 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_585
timestamp 1644511149
transform 1 0 54924 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_597
timestamp 1644511149
transform 1 0 56028 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_609
timestamp 1644511149
transform 1 0 57132 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_615
timestamp 1644511149
transform 1 0 57684 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_43_617
timestamp 1644511149
transform 1 0 57868 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_44_3
timestamp 1644511149
transform 1 0 1380 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_15
timestamp 1644511149
transform 1 0 2484 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_44_27
timestamp 1644511149
transform 1 0 3588 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_29
timestamp 1644511149
transform 1 0 3772 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_41
timestamp 1644511149
transform 1 0 4876 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_53
timestamp 1644511149
transform 1 0 5980 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_65
timestamp 1644511149
transform 1 0 7084 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_77
timestamp 1644511149
transform 1 0 8188 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_83
timestamp 1644511149
transform 1 0 8740 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_85
timestamp 1644511149
transform 1 0 8924 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_97
timestamp 1644511149
transform 1 0 10028 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_109
timestamp 1644511149
transform 1 0 11132 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_121
timestamp 1644511149
transform 1 0 12236 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_133
timestamp 1644511149
transform 1 0 13340 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_139
timestamp 1644511149
transform 1 0 13892 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_141
timestamp 1644511149
transform 1 0 14076 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_153
timestamp 1644511149
transform 1 0 15180 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_165
timestamp 1644511149
transform 1 0 16284 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_177
timestamp 1644511149
transform 1 0 17388 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_189
timestamp 1644511149
transform 1 0 18492 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_195
timestamp 1644511149
transform 1 0 19044 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_197
timestamp 1644511149
transform 1 0 19228 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_209
timestamp 1644511149
transform 1 0 20332 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_221
timestamp 1644511149
transform 1 0 21436 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_233
timestamp 1644511149
transform 1 0 22540 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_245
timestamp 1644511149
transform 1 0 23644 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_251
timestamp 1644511149
transform 1 0 24196 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_253
timestamp 1644511149
transform 1 0 24380 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_265
timestamp 1644511149
transform 1 0 25484 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_277
timestamp 1644511149
transform 1 0 26588 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_289
timestamp 1644511149
transform 1 0 27692 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_301
timestamp 1644511149
transform 1 0 28796 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_307
timestamp 1644511149
transform 1 0 29348 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_309
timestamp 1644511149
transform 1 0 29532 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_321
timestamp 1644511149
transform 1 0 30636 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_333
timestamp 1644511149
transform 1 0 31740 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_345
timestamp 1644511149
transform 1 0 32844 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_357
timestamp 1644511149
transform 1 0 33948 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_363
timestamp 1644511149
transform 1 0 34500 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_365
timestamp 1644511149
transform 1 0 34684 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_377
timestamp 1644511149
transform 1 0 35788 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_389
timestamp 1644511149
transform 1 0 36892 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_401
timestamp 1644511149
transform 1 0 37996 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_413
timestamp 1644511149
transform 1 0 39100 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_419
timestamp 1644511149
transform 1 0 39652 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_421
timestamp 1644511149
transform 1 0 39836 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_433
timestamp 1644511149
transform 1 0 40940 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_445
timestamp 1644511149
transform 1 0 42044 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_457
timestamp 1644511149
transform 1 0 43148 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_469
timestamp 1644511149
transform 1 0 44252 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_475
timestamp 1644511149
transform 1 0 44804 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_477
timestamp 1644511149
transform 1 0 44988 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_489
timestamp 1644511149
transform 1 0 46092 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_501
timestamp 1644511149
transform 1 0 47196 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_513
timestamp 1644511149
transform 1 0 48300 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_525
timestamp 1644511149
transform 1 0 49404 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_531
timestamp 1644511149
transform 1 0 49956 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_533
timestamp 1644511149
transform 1 0 50140 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_545
timestamp 1644511149
transform 1 0 51244 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_557
timestamp 1644511149
transform 1 0 52348 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_569
timestamp 1644511149
transform 1 0 53452 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_581
timestamp 1644511149
transform 1 0 54556 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_587
timestamp 1644511149
transform 1 0 55108 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_589
timestamp 1644511149
transform 1 0 55292 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_601
timestamp 1644511149
transform 1 0 56396 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_613
timestamp 1644511149
transform 1 0 57500 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_3
timestamp 1644511149
transform 1 0 1380 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_15
timestamp 1644511149
transform 1 0 2484 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_27
timestamp 1644511149
transform 1 0 3588 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_39
timestamp 1644511149
transform 1 0 4692 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_51
timestamp 1644511149
transform 1 0 5796 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_55
timestamp 1644511149
transform 1 0 6164 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_57
timestamp 1644511149
transform 1 0 6348 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_69
timestamp 1644511149
transform 1 0 7452 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_81
timestamp 1644511149
transform 1 0 8556 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_93
timestamp 1644511149
transform 1 0 9660 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_105
timestamp 1644511149
transform 1 0 10764 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_111
timestamp 1644511149
transform 1 0 11316 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_113
timestamp 1644511149
transform 1 0 11500 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_125
timestamp 1644511149
transform 1 0 12604 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_137
timestamp 1644511149
transform 1 0 13708 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_149
timestamp 1644511149
transform 1 0 14812 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_161
timestamp 1644511149
transform 1 0 15916 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_167
timestamp 1644511149
transform 1 0 16468 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_169
timestamp 1644511149
transform 1 0 16652 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_181
timestamp 1644511149
transform 1 0 17756 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_193
timestamp 1644511149
transform 1 0 18860 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_205
timestamp 1644511149
transform 1 0 19964 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_217
timestamp 1644511149
transform 1 0 21068 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_223
timestamp 1644511149
transform 1 0 21620 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_225
timestamp 1644511149
transform 1 0 21804 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_237
timestamp 1644511149
transform 1 0 22908 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_249
timestamp 1644511149
transform 1 0 24012 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_261
timestamp 1644511149
transform 1 0 25116 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_273
timestamp 1644511149
transform 1 0 26220 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_279
timestamp 1644511149
transform 1 0 26772 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_281
timestamp 1644511149
transform 1 0 26956 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_293
timestamp 1644511149
transform 1 0 28060 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_305
timestamp 1644511149
transform 1 0 29164 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_317
timestamp 1644511149
transform 1 0 30268 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_329
timestamp 1644511149
transform 1 0 31372 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_335
timestamp 1644511149
transform 1 0 31924 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_337
timestamp 1644511149
transform 1 0 32108 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_349
timestamp 1644511149
transform 1 0 33212 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_361
timestamp 1644511149
transform 1 0 34316 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_373
timestamp 1644511149
transform 1 0 35420 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_385
timestamp 1644511149
transform 1 0 36524 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_391
timestamp 1644511149
transform 1 0 37076 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_393
timestamp 1644511149
transform 1 0 37260 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_405
timestamp 1644511149
transform 1 0 38364 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_417
timestamp 1644511149
transform 1 0 39468 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_429
timestamp 1644511149
transform 1 0 40572 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_441
timestamp 1644511149
transform 1 0 41676 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_447
timestamp 1644511149
transform 1 0 42228 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_449
timestamp 1644511149
transform 1 0 42412 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_461
timestamp 1644511149
transform 1 0 43516 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_473
timestamp 1644511149
transform 1 0 44620 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_485
timestamp 1644511149
transform 1 0 45724 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_497
timestamp 1644511149
transform 1 0 46828 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_503
timestamp 1644511149
transform 1 0 47380 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_505
timestamp 1644511149
transform 1 0 47564 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_517
timestamp 1644511149
transform 1 0 48668 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_529
timestamp 1644511149
transform 1 0 49772 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_541
timestamp 1644511149
transform 1 0 50876 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_553
timestamp 1644511149
transform 1 0 51980 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_559
timestamp 1644511149
transform 1 0 52532 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_561
timestamp 1644511149
transform 1 0 52716 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_573
timestamp 1644511149
transform 1 0 53820 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_585
timestamp 1644511149
transform 1 0 54924 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_597
timestamp 1644511149
transform 1 0 56028 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_609
timestamp 1644511149
transform 1 0 57132 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_615
timestamp 1644511149
transform 1 0 57684 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_45_617
timestamp 1644511149
transform 1 0 57868 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_46_3
timestamp 1644511149
transform 1 0 1380 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_15
timestamp 1644511149
transform 1 0 2484 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_46_27
timestamp 1644511149
transform 1 0 3588 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_29
timestamp 1644511149
transform 1 0 3772 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_41
timestamp 1644511149
transform 1 0 4876 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_53
timestamp 1644511149
transform 1 0 5980 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_65
timestamp 1644511149
transform 1 0 7084 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_77
timestamp 1644511149
transform 1 0 8188 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_83
timestamp 1644511149
transform 1 0 8740 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_85
timestamp 1644511149
transform 1 0 8924 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_97
timestamp 1644511149
transform 1 0 10028 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_109
timestamp 1644511149
transform 1 0 11132 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_121
timestamp 1644511149
transform 1 0 12236 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_133
timestamp 1644511149
transform 1 0 13340 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_139
timestamp 1644511149
transform 1 0 13892 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_141
timestamp 1644511149
transform 1 0 14076 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_153
timestamp 1644511149
transform 1 0 15180 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_165
timestamp 1644511149
transform 1 0 16284 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_177
timestamp 1644511149
transform 1 0 17388 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_189
timestamp 1644511149
transform 1 0 18492 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_195
timestamp 1644511149
transform 1 0 19044 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_197
timestamp 1644511149
transform 1 0 19228 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_209
timestamp 1644511149
transform 1 0 20332 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_221
timestamp 1644511149
transform 1 0 21436 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_233
timestamp 1644511149
transform 1 0 22540 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_245
timestamp 1644511149
transform 1 0 23644 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_251
timestamp 1644511149
transform 1 0 24196 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_253
timestamp 1644511149
transform 1 0 24380 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_265
timestamp 1644511149
transform 1 0 25484 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_277
timestamp 1644511149
transform 1 0 26588 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_289
timestamp 1644511149
transform 1 0 27692 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_301
timestamp 1644511149
transform 1 0 28796 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_307
timestamp 1644511149
transform 1 0 29348 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_309
timestamp 1644511149
transform 1 0 29532 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_321
timestamp 1644511149
transform 1 0 30636 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_333
timestamp 1644511149
transform 1 0 31740 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_345
timestamp 1644511149
transform 1 0 32844 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_357
timestamp 1644511149
transform 1 0 33948 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_363
timestamp 1644511149
transform 1 0 34500 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_365
timestamp 1644511149
transform 1 0 34684 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_377
timestamp 1644511149
transform 1 0 35788 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_389
timestamp 1644511149
transform 1 0 36892 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_401
timestamp 1644511149
transform 1 0 37996 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_413
timestamp 1644511149
transform 1 0 39100 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_419
timestamp 1644511149
transform 1 0 39652 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_421
timestamp 1644511149
transform 1 0 39836 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_433
timestamp 1644511149
transform 1 0 40940 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_445
timestamp 1644511149
transform 1 0 42044 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_457
timestamp 1644511149
transform 1 0 43148 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_469
timestamp 1644511149
transform 1 0 44252 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_475
timestamp 1644511149
transform 1 0 44804 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_477
timestamp 1644511149
transform 1 0 44988 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_489
timestamp 1644511149
transform 1 0 46092 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_501
timestamp 1644511149
transform 1 0 47196 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_513
timestamp 1644511149
transform 1 0 48300 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_525
timestamp 1644511149
transform 1 0 49404 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_531
timestamp 1644511149
transform 1 0 49956 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_533
timestamp 1644511149
transform 1 0 50140 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_545
timestamp 1644511149
transform 1 0 51244 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_557
timestamp 1644511149
transform 1 0 52348 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_569
timestamp 1644511149
transform 1 0 53452 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_581
timestamp 1644511149
transform 1 0 54556 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_587
timestamp 1644511149
transform 1 0 55108 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_589
timestamp 1644511149
transform 1 0 55292 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_601
timestamp 1644511149
transform 1 0 56396 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_613
timestamp 1644511149
transform 1 0 57500 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_3
timestamp 1644511149
transform 1 0 1380 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_15
timestamp 1644511149
transform 1 0 2484 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_27
timestamp 1644511149
transform 1 0 3588 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_39
timestamp 1644511149
transform 1 0 4692 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_51
timestamp 1644511149
transform 1 0 5796 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_55
timestamp 1644511149
transform 1 0 6164 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_57
timestamp 1644511149
transform 1 0 6348 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_69
timestamp 1644511149
transform 1 0 7452 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_81
timestamp 1644511149
transform 1 0 8556 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_93
timestamp 1644511149
transform 1 0 9660 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_105
timestamp 1644511149
transform 1 0 10764 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_111
timestamp 1644511149
transform 1 0 11316 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_113
timestamp 1644511149
transform 1 0 11500 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_125
timestamp 1644511149
transform 1 0 12604 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_137
timestamp 1644511149
transform 1 0 13708 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_149
timestamp 1644511149
transform 1 0 14812 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_161
timestamp 1644511149
transform 1 0 15916 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_167
timestamp 1644511149
transform 1 0 16468 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_169
timestamp 1644511149
transform 1 0 16652 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_181
timestamp 1644511149
transform 1 0 17756 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_193
timestamp 1644511149
transform 1 0 18860 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_205
timestamp 1644511149
transform 1 0 19964 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_217
timestamp 1644511149
transform 1 0 21068 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_223
timestamp 1644511149
transform 1 0 21620 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_225
timestamp 1644511149
transform 1 0 21804 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_237
timestamp 1644511149
transform 1 0 22908 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_249
timestamp 1644511149
transform 1 0 24012 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_261
timestamp 1644511149
transform 1 0 25116 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_273
timestamp 1644511149
transform 1 0 26220 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_279
timestamp 1644511149
transform 1 0 26772 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_281
timestamp 1644511149
transform 1 0 26956 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_293
timestamp 1644511149
transform 1 0 28060 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_305
timestamp 1644511149
transform 1 0 29164 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_317
timestamp 1644511149
transform 1 0 30268 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_329
timestamp 1644511149
transform 1 0 31372 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_335
timestamp 1644511149
transform 1 0 31924 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_337
timestamp 1644511149
transform 1 0 32108 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_349
timestamp 1644511149
transform 1 0 33212 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_361
timestamp 1644511149
transform 1 0 34316 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_373
timestamp 1644511149
transform 1 0 35420 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_385
timestamp 1644511149
transform 1 0 36524 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_391
timestamp 1644511149
transform 1 0 37076 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_393
timestamp 1644511149
transform 1 0 37260 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_405
timestamp 1644511149
transform 1 0 38364 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_417
timestamp 1644511149
transform 1 0 39468 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_429
timestamp 1644511149
transform 1 0 40572 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_441
timestamp 1644511149
transform 1 0 41676 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_447
timestamp 1644511149
transform 1 0 42228 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_449
timestamp 1644511149
transform 1 0 42412 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_461
timestamp 1644511149
transform 1 0 43516 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_473
timestamp 1644511149
transform 1 0 44620 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_485
timestamp 1644511149
transform 1 0 45724 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_497
timestamp 1644511149
transform 1 0 46828 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_503
timestamp 1644511149
transform 1 0 47380 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_505
timestamp 1644511149
transform 1 0 47564 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_517
timestamp 1644511149
transform 1 0 48668 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_529
timestamp 1644511149
transform 1 0 49772 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_541
timestamp 1644511149
transform 1 0 50876 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_553
timestamp 1644511149
transform 1 0 51980 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_559
timestamp 1644511149
transform 1 0 52532 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_561
timestamp 1644511149
transform 1 0 52716 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_573
timestamp 1644511149
transform 1 0 53820 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_585
timestamp 1644511149
transform 1 0 54924 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_597
timestamp 1644511149
transform 1 0 56028 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_609
timestamp 1644511149
transform 1 0 57132 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_615
timestamp 1644511149
transform 1 0 57684 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_47_617
timestamp 1644511149
transform 1 0 57868 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_48_3
timestamp 1644511149
transform 1 0 1380 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_15
timestamp 1644511149
transform 1 0 2484 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_48_27
timestamp 1644511149
transform 1 0 3588 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_29
timestamp 1644511149
transform 1 0 3772 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_41
timestamp 1644511149
transform 1 0 4876 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_53
timestamp 1644511149
transform 1 0 5980 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_65
timestamp 1644511149
transform 1 0 7084 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_77
timestamp 1644511149
transform 1 0 8188 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_83
timestamp 1644511149
transform 1 0 8740 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_85
timestamp 1644511149
transform 1 0 8924 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_97
timestamp 1644511149
transform 1 0 10028 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_109
timestamp 1644511149
transform 1 0 11132 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_121
timestamp 1644511149
transform 1 0 12236 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_133
timestamp 1644511149
transform 1 0 13340 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_139
timestamp 1644511149
transform 1 0 13892 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_141
timestamp 1644511149
transform 1 0 14076 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_153
timestamp 1644511149
transform 1 0 15180 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_165
timestamp 1644511149
transform 1 0 16284 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_177
timestamp 1644511149
transform 1 0 17388 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_189
timestamp 1644511149
transform 1 0 18492 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_195
timestamp 1644511149
transform 1 0 19044 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_197
timestamp 1644511149
transform 1 0 19228 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_209
timestamp 1644511149
transform 1 0 20332 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_221
timestamp 1644511149
transform 1 0 21436 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_233
timestamp 1644511149
transform 1 0 22540 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_245
timestamp 1644511149
transform 1 0 23644 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_251
timestamp 1644511149
transform 1 0 24196 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_253
timestamp 1644511149
transform 1 0 24380 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_265
timestamp 1644511149
transform 1 0 25484 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_277
timestamp 1644511149
transform 1 0 26588 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_289
timestamp 1644511149
transform 1 0 27692 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_301
timestamp 1644511149
transform 1 0 28796 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_307
timestamp 1644511149
transform 1 0 29348 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_309
timestamp 1644511149
transform 1 0 29532 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_321
timestamp 1644511149
transform 1 0 30636 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_333
timestamp 1644511149
transform 1 0 31740 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_345
timestamp 1644511149
transform 1 0 32844 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_357
timestamp 1644511149
transform 1 0 33948 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_363
timestamp 1644511149
transform 1 0 34500 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_365
timestamp 1644511149
transform 1 0 34684 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_377
timestamp 1644511149
transform 1 0 35788 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_389
timestamp 1644511149
transform 1 0 36892 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_401
timestamp 1644511149
transform 1 0 37996 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_413
timestamp 1644511149
transform 1 0 39100 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_419
timestamp 1644511149
transform 1 0 39652 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_421
timestamp 1644511149
transform 1 0 39836 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_433
timestamp 1644511149
transform 1 0 40940 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_445
timestamp 1644511149
transform 1 0 42044 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_457
timestamp 1644511149
transform 1 0 43148 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_469
timestamp 1644511149
transform 1 0 44252 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_475
timestamp 1644511149
transform 1 0 44804 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_477
timestamp 1644511149
transform 1 0 44988 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_489
timestamp 1644511149
transform 1 0 46092 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_501
timestamp 1644511149
transform 1 0 47196 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_513
timestamp 1644511149
transform 1 0 48300 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_525
timestamp 1644511149
transform 1 0 49404 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_531
timestamp 1644511149
transform 1 0 49956 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_533
timestamp 1644511149
transform 1 0 50140 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_545
timestamp 1644511149
transform 1 0 51244 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_557
timestamp 1644511149
transform 1 0 52348 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_569
timestamp 1644511149
transform 1 0 53452 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_581
timestamp 1644511149
transform 1 0 54556 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_587
timestamp 1644511149
transform 1 0 55108 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_48_589
timestamp 1644511149
transform 1 0 55292 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_48_597
timestamp 1644511149
transform 1 0 56028 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_48_621
timestamp 1644511149
transform 1 0 58236 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_49_3
timestamp 1644511149
transform 1 0 1380 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_15
timestamp 1644511149
transform 1 0 2484 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_27
timestamp 1644511149
transform 1 0 3588 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_39
timestamp 1644511149
transform 1 0 4692 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_51
timestamp 1644511149
transform 1 0 5796 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_55
timestamp 1644511149
transform 1 0 6164 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_57
timestamp 1644511149
transform 1 0 6348 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_69
timestamp 1644511149
transform 1 0 7452 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_81
timestamp 1644511149
transform 1 0 8556 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_93
timestamp 1644511149
transform 1 0 9660 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_105
timestamp 1644511149
transform 1 0 10764 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_111
timestamp 1644511149
transform 1 0 11316 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_113
timestamp 1644511149
transform 1 0 11500 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_125
timestamp 1644511149
transform 1 0 12604 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_137
timestamp 1644511149
transform 1 0 13708 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_149
timestamp 1644511149
transform 1 0 14812 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_161
timestamp 1644511149
transform 1 0 15916 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_167
timestamp 1644511149
transform 1 0 16468 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_169
timestamp 1644511149
transform 1 0 16652 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_181
timestamp 1644511149
transform 1 0 17756 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_193
timestamp 1644511149
transform 1 0 18860 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_205
timestamp 1644511149
transform 1 0 19964 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_217
timestamp 1644511149
transform 1 0 21068 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_223
timestamp 1644511149
transform 1 0 21620 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_225
timestamp 1644511149
transform 1 0 21804 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_237
timestamp 1644511149
transform 1 0 22908 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_249
timestamp 1644511149
transform 1 0 24012 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_261
timestamp 1644511149
transform 1 0 25116 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_273
timestamp 1644511149
transform 1 0 26220 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_279
timestamp 1644511149
transform 1 0 26772 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_281
timestamp 1644511149
transform 1 0 26956 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_293
timestamp 1644511149
transform 1 0 28060 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_305
timestamp 1644511149
transform 1 0 29164 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_317
timestamp 1644511149
transform 1 0 30268 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_329
timestamp 1644511149
transform 1 0 31372 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_335
timestamp 1644511149
transform 1 0 31924 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_337
timestamp 1644511149
transform 1 0 32108 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_349
timestamp 1644511149
transform 1 0 33212 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_361
timestamp 1644511149
transform 1 0 34316 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_373
timestamp 1644511149
transform 1 0 35420 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_385
timestamp 1644511149
transform 1 0 36524 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_391
timestamp 1644511149
transform 1 0 37076 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_393
timestamp 1644511149
transform 1 0 37260 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_405
timestamp 1644511149
transform 1 0 38364 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_417
timestamp 1644511149
transform 1 0 39468 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_429
timestamp 1644511149
transform 1 0 40572 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_441
timestamp 1644511149
transform 1 0 41676 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_447
timestamp 1644511149
transform 1 0 42228 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_449
timestamp 1644511149
transform 1 0 42412 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_461
timestamp 1644511149
transform 1 0 43516 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_473
timestamp 1644511149
transform 1 0 44620 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_485
timestamp 1644511149
transform 1 0 45724 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_497
timestamp 1644511149
transform 1 0 46828 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_503
timestamp 1644511149
transform 1 0 47380 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_505
timestamp 1644511149
transform 1 0 47564 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_517
timestamp 1644511149
transform 1 0 48668 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_529
timestamp 1644511149
transform 1 0 49772 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_541
timestamp 1644511149
transform 1 0 50876 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_553
timestamp 1644511149
transform 1 0 51980 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_559
timestamp 1644511149
transform 1 0 52532 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_561
timestamp 1644511149
transform 1 0 52716 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_573
timestamp 1644511149
transform 1 0 53820 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_585
timestamp 1644511149
transform 1 0 54924 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_49_597
timestamp 1644511149
transform 1 0 56028 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_49_605
timestamp 1644511149
transform 1 0 56764 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_49_610
timestamp 1644511149
transform 1 0 57224 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_49_620
timestamp 1644511149
transform 1 0 58144 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_624
timestamp 1644511149
transform 1 0 58512 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_3
timestamp 1644511149
transform 1 0 1380 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_15
timestamp 1644511149
transform 1 0 2484 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_50_27
timestamp 1644511149
transform 1 0 3588 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_29
timestamp 1644511149
transform 1 0 3772 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_41
timestamp 1644511149
transform 1 0 4876 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_53
timestamp 1644511149
transform 1 0 5980 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_65
timestamp 1644511149
transform 1 0 7084 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_77
timestamp 1644511149
transform 1 0 8188 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_83
timestamp 1644511149
transform 1 0 8740 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_85
timestamp 1644511149
transform 1 0 8924 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_97
timestamp 1644511149
transform 1 0 10028 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_109
timestamp 1644511149
transform 1 0 11132 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_121
timestamp 1644511149
transform 1 0 12236 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_133
timestamp 1644511149
transform 1 0 13340 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_139
timestamp 1644511149
transform 1 0 13892 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_141
timestamp 1644511149
transform 1 0 14076 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_153
timestamp 1644511149
transform 1 0 15180 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_165
timestamp 1644511149
transform 1 0 16284 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_177
timestamp 1644511149
transform 1 0 17388 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_189
timestamp 1644511149
transform 1 0 18492 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_195
timestamp 1644511149
transform 1 0 19044 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_197
timestamp 1644511149
transform 1 0 19228 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_209
timestamp 1644511149
transform 1 0 20332 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_221
timestamp 1644511149
transform 1 0 21436 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_233
timestamp 1644511149
transform 1 0 22540 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_245
timestamp 1644511149
transform 1 0 23644 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_251
timestamp 1644511149
transform 1 0 24196 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_253
timestamp 1644511149
transform 1 0 24380 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_265
timestamp 1644511149
transform 1 0 25484 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_277
timestamp 1644511149
transform 1 0 26588 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_289
timestamp 1644511149
transform 1 0 27692 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_301
timestamp 1644511149
transform 1 0 28796 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_307
timestamp 1644511149
transform 1 0 29348 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_309
timestamp 1644511149
transform 1 0 29532 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_321
timestamp 1644511149
transform 1 0 30636 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_333
timestamp 1644511149
transform 1 0 31740 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_345
timestamp 1644511149
transform 1 0 32844 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_357
timestamp 1644511149
transform 1 0 33948 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_363
timestamp 1644511149
transform 1 0 34500 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_365
timestamp 1644511149
transform 1 0 34684 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_377
timestamp 1644511149
transform 1 0 35788 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_389
timestamp 1644511149
transform 1 0 36892 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_401
timestamp 1644511149
transform 1 0 37996 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_413
timestamp 1644511149
transform 1 0 39100 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_419
timestamp 1644511149
transform 1 0 39652 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_421
timestamp 1644511149
transform 1 0 39836 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_433
timestamp 1644511149
transform 1 0 40940 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_445
timestamp 1644511149
transform 1 0 42044 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_457
timestamp 1644511149
transform 1 0 43148 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_469
timestamp 1644511149
transform 1 0 44252 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_475
timestamp 1644511149
transform 1 0 44804 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_477
timestamp 1644511149
transform 1 0 44988 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_489
timestamp 1644511149
transform 1 0 46092 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_501
timestamp 1644511149
transform 1 0 47196 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_513
timestamp 1644511149
transform 1 0 48300 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_525
timestamp 1644511149
transform 1 0 49404 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_531
timestamp 1644511149
transform 1 0 49956 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_533
timestamp 1644511149
transform 1 0 50140 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_545
timestamp 1644511149
transform 1 0 51244 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_557
timestamp 1644511149
transform 1 0 52348 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_569
timestamp 1644511149
transform 1 0 53452 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_581
timestamp 1644511149
transform 1 0 54556 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_587
timestamp 1644511149
transform 1 0 55108 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_589
timestamp 1644511149
transform 1 0 55292 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_601
timestamp 1644511149
transform 1 0 56396 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_613
timestamp 1644511149
transform 1 0 57500 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_3
timestamp 1644511149
transform 1 0 1380 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_15
timestamp 1644511149
transform 1 0 2484 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_27
timestamp 1644511149
transform 1 0 3588 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_39
timestamp 1644511149
transform 1 0 4692 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_51
timestamp 1644511149
transform 1 0 5796 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_55
timestamp 1644511149
transform 1 0 6164 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_57
timestamp 1644511149
transform 1 0 6348 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_69
timestamp 1644511149
transform 1 0 7452 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_81
timestamp 1644511149
transform 1 0 8556 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_93
timestamp 1644511149
transform 1 0 9660 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_105
timestamp 1644511149
transform 1 0 10764 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_111
timestamp 1644511149
transform 1 0 11316 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_113
timestamp 1644511149
transform 1 0 11500 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_125
timestamp 1644511149
transform 1 0 12604 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_137
timestamp 1644511149
transform 1 0 13708 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_149
timestamp 1644511149
transform 1 0 14812 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_161
timestamp 1644511149
transform 1 0 15916 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_167
timestamp 1644511149
transform 1 0 16468 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_169
timestamp 1644511149
transform 1 0 16652 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_181
timestamp 1644511149
transform 1 0 17756 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_193
timestamp 1644511149
transform 1 0 18860 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_205
timestamp 1644511149
transform 1 0 19964 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_217
timestamp 1644511149
transform 1 0 21068 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_223
timestamp 1644511149
transform 1 0 21620 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_225
timestamp 1644511149
transform 1 0 21804 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_237
timestamp 1644511149
transform 1 0 22908 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_249
timestamp 1644511149
transform 1 0 24012 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_261
timestamp 1644511149
transform 1 0 25116 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_273
timestamp 1644511149
transform 1 0 26220 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_279
timestamp 1644511149
transform 1 0 26772 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_281
timestamp 1644511149
transform 1 0 26956 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_293
timestamp 1644511149
transform 1 0 28060 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_305
timestamp 1644511149
transform 1 0 29164 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_317
timestamp 1644511149
transform 1 0 30268 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_329
timestamp 1644511149
transform 1 0 31372 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_335
timestamp 1644511149
transform 1 0 31924 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_337
timestamp 1644511149
transform 1 0 32108 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_349
timestamp 1644511149
transform 1 0 33212 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_361
timestamp 1644511149
transform 1 0 34316 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_373
timestamp 1644511149
transform 1 0 35420 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_385
timestamp 1644511149
transform 1 0 36524 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_391
timestamp 1644511149
transform 1 0 37076 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_393
timestamp 1644511149
transform 1 0 37260 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_405
timestamp 1644511149
transform 1 0 38364 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_417
timestamp 1644511149
transform 1 0 39468 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_429
timestamp 1644511149
transform 1 0 40572 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_441
timestamp 1644511149
transform 1 0 41676 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_447
timestamp 1644511149
transform 1 0 42228 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_449
timestamp 1644511149
transform 1 0 42412 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_461
timestamp 1644511149
transform 1 0 43516 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_473
timestamp 1644511149
transform 1 0 44620 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_485
timestamp 1644511149
transform 1 0 45724 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_497
timestamp 1644511149
transform 1 0 46828 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_503
timestamp 1644511149
transform 1 0 47380 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_505
timestamp 1644511149
transform 1 0 47564 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_517
timestamp 1644511149
transform 1 0 48668 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_529
timestamp 1644511149
transform 1 0 49772 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_541
timestamp 1644511149
transform 1 0 50876 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_553
timestamp 1644511149
transform 1 0 51980 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_559
timestamp 1644511149
transform 1 0 52532 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_561
timestamp 1644511149
transform 1 0 52716 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_573
timestamp 1644511149
transform 1 0 53820 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_585
timestamp 1644511149
transform 1 0 54924 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_597
timestamp 1644511149
transform 1 0 56028 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_609
timestamp 1644511149
transform 1 0 57132 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_615
timestamp 1644511149
transform 1 0 57684 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_51_617
timestamp 1644511149
transform 1 0 57868 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_52_3
timestamp 1644511149
transform 1 0 1380 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_15
timestamp 1644511149
transform 1 0 2484 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_52_27
timestamp 1644511149
transform 1 0 3588 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_29
timestamp 1644511149
transform 1 0 3772 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_41
timestamp 1644511149
transform 1 0 4876 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_53
timestamp 1644511149
transform 1 0 5980 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_65
timestamp 1644511149
transform 1 0 7084 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_77
timestamp 1644511149
transform 1 0 8188 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_83
timestamp 1644511149
transform 1 0 8740 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_85
timestamp 1644511149
transform 1 0 8924 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_97
timestamp 1644511149
transform 1 0 10028 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_109
timestamp 1644511149
transform 1 0 11132 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_121
timestamp 1644511149
transform 1 0 12236 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_133
timestamp 1644511149
transform 1 0 13340 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_139
timestamp 1644511149
transform 1 0 13892 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_141
timestamp 1644511149
transform 1 0 14076 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_153
timestamp 1644511149
transform 1 0 15180 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_165
timestamp 1644511149
transform 1 0 16284 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_177
timestamp 1644511149
transform 1 0 17388 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_189
timestamp 1644511149
transform 1 0 18492 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_195
timestamp 1644511149
transform 1 0 19044 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_197
timestamp 1644511149
transform 1 0 19228 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_209
timestamp 1644511149
transform 1 0 20332 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_221
timestamp 1644511149
transform 1 0 21436 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_233
timestamp 1644511149
transform 1 0 22540 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_245
timestamp 1644511149
transform 1 0 23644 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_251
timestamp 1644511149
transform 1 0 24196 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_253
timestamp 1644511149
transform 1 0 24380 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_265
timestamp 1644511149
transform 1 0 25484 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_277
timestamp 1644511149
transform 1 0 26588 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_289
timestamp 1644511149
transform 1 0 27692 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_301
timestamp 1644511149
transform 1 0 28796 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_307
timestamp 1644511149
transform 1 0 29348 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_309
timestamp 1644511149
transform 1 0 29532 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_321
timestamp 1644511149
transform 1 0 30636 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_333
timestamp 1644511149
transform 1 0 31740 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_345
timestamp 1644511149
transform 1 0 32844 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_357
timestamp 1644511149
transform 1 0 33948 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_363
timestamp 1644511149
transform 1 0 34500 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_365
timestamp 1644511149
transform 1 0 34684 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_377
timestamp 1644511149
transform 1 0 35788 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_389
timestamp 1644511149
transform 1 0 36892 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_401
timestamp 1644511149
transform 1 0 37996 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_413
timestamp 1644511149
transform 1 0 39100 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_419
timestamp 1644511149
transform 1 0 39652 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_421
timestamp 1644511149
transform 1 0 39836 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_433
timestamp 1644511149
transform 1 0 40940 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_445
timestamp 1644511149
transform 1 0 42044 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_457
timestamp 1644511149
transform 1 0 43148 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_469
timestamp 1644511149
transform 1 0 44252 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_475
timestamp 1644511149
transform 1 0 44804 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_477
timestamp 1644511149
transform 1 0 44988 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_489
timestamp 1644511149
transform 1 0 46092 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_501
timestamp 1644511149
transform 1 0 47196 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_513
timestamp 1644511149
transform 1 0 48300 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_525
timestamp 1644511149
transform 1 0 49404 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_531
timestamp 1644511149
transform 1 0 49956 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_533
timestamp 1644511149
transform 1 0 50140 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_545
timestamp 1644511149
transform 1 0 51244 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_557
timestamp 1644511149
transform 1 0 52348 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_569
timestamp 1644511149
transform 1 0 53452 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_581
timestamp 1644511149
transform 1 0 54556 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_587
timestamp 1644511149
transform 1 0 55108 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_589
timestamp 1644511149
transform 1 0 55292 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_601
timestamp 1644511149
transform 1 0 56396 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_613
timestamp 1644511149
transform 1 0 57500 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_3
timestamp 1644511149
transform 1 0 1380 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_15
timestamp 1644511149
transform 1 0 2484 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_27
timestamp 1644511149
transform 1 0 3588 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_39
timestamp 1644511149
transform 1 0 4692 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_51
timestamp 1644511149
transform 1 0 5796 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_55
timestamp 1644511149
transform 1 0 6164 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_57
timestamp 1644511149
transform 1 0 6348 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_69
timestamp 1644511149
transform 1 0 7452 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_81
timestamp 1644511149
transform 1 0 8556 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_93
timestamp 1644511149
transform 1 0 9660 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_105
timestamp 1644511149
transform 1 0 10764 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_111
timestamp 1644511149
transform 1 0 11316 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_113
timestamp 1644511149
transform 1 0 11500 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_125
timestamp 1644511149
transform 1 0 12604 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_137
timestamp 1644511149
transform 1 0 13708 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_149
timestamp 1644511149
transform 1 0 14812 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_161
timestamp 1644511149
transform 1 0 15916 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_167
timestamp 1644511149
transform 1 0 16468 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_169
timestamp 1644511149
transform 1 0 16652 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_181
timestamp 1644511149
transform 1 0 17756 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_193
timestamp 1644511149
transform 1 0 18860 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_205
timestamp 1644511149
transform 1 0 19964 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_217
timestamp 1644511149
transform 1 0 21068 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_223
timestamp 1644511149
transform 1 0 21620 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_225
timestamp 1644511149
transform 1 0 21804 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_237
timestamp 1644511149
transform 1 0 22908 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_249
timestamp 1644511149
transform 1 0 24012 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_261
timestamp 1644511149
transform 1 0 25116 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_273
timestamp 1644511149
transform 1 0 26220 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_279
timestamp 1644511149
transform 1 0 26772 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_281
timestamp 1644511149
transform 1 0 26956 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_293
timestamp 1644511149
transform 1 0 28060 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_305
timestamp 1644511149
transform 1 0 29164 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_317
timestamp 1644511149
transform 1 0 30268 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_329
timestamp 1644511149
transform 1 0 31372 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_335
timestamp 1644511149
transform 1 0 31924 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_337
timestamp 1644511149
transform 1 0 32108 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_349
timestamp 1644511149
transform 1 0 33212 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_361
timestamp 1644511149
transform 1 0 34316 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_373
timestamp 1644511149
transform 1 0 35420 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_385
timestamp 1644511149
transform 1 0 36524 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_391
timestamp 1644511149
transform 1 0 37076 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_393
timestamp 1644511149
transform 1 0 37260 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_405
timestamp 1644511149
transform 1 0 38364 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_417
timestamp 1644511149
transform 1 0 39468 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_429
timestamp 1644511149
transform 1 0 40572 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_441
timestamp 1644511149
transform 1 0 41676 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_447
timestamp 1644511149
transform 1 0 42228 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_449
timestamp 1644511149
transform 1 0 42412 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_461
timestamp 1644511149
transform 1 0 43516 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_473
timestamp 1644511149
transform 1 0 44620 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_485
timestamp 1644511149
transform 1 0 45724 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_497
timestamp 1644511149
transform 1 0 46828 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_503
timestamp 1644511149
transform 1 0 47380 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_505
timestamp 1644511149
transform 1 0 47564 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_517
timestamp 1644511149
transform 1 0 48668 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_529
timestamp 1644511149
transform 1 0 49772 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_541
timestamp 1644511149
transform 1 0 50876 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_553
timestamp 1644511149
transform 1 0 51980 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_559
timestamp 1644511149
transform 1 0 52532 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_561
timestamp 1644511149
transform 1 0 52716 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_573
timestamp 1644511149
transform 1 0 53820 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_585
timestamp 1644511149
transform 1 0 54924 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_597
timestamp 1644511149
transform 1 0 56028 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_609
timestamp 1644511149
transform 1 0 57132 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_615
timestamp 1644511149
transform 1 0 57684 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_53_617
timestamp 1644511149
transform 1 0 57868 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_54_3
timestamp 1644511149
transform 1 0 1380 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_15
timestamp 1644511149
transform 1 0 2484 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_54_27
timestamp 1644511149
transform 1 0 3588 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_29
timestamp 1644511149
transform 1 0 3772 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_41
timestamp 1644511149
transform 1 0 4876 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_53
timestamp 1644511149
transform 1 0 5980 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_65
timestamp 1644511149
transform 1 0 7084 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_77
timestamp 1644511149
transform 1 0 8188 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_83
timestamp 1644511149
transform 1 0 8740 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_85
timestamp 1644511149
transform 1 0 8924 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_97
timestamp 1644511149
transform 1 0 10028 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_109
timestamp 1644511149
transform 1 0 11132 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_121
timestamp 1644511149
transform 1 0 12236 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_133
timestamp 1644511149
transform 1 0 13340 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_139
timestamp 1644511149
transform 1 0 13892 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_141
timestamp 1644511149
transform 1 0 14076 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_153
timestamp 1644511149
transform 1 0 15180 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_165
timestamp 1644511149
transform 1 0 16284 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_177
timestamp 1644511149
transform 1 0 17388 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_189
timestamp 1644511149
transform 1 0 18492 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_195
timestamp 1644511149
transform 1 0 19044 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_197
timestamp 1644511149
transform 1 0 19228 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_209
timestamp 1644511149
transform 1 0 20332 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_221
timestamp 1644511149
transform 1 0 21436 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_233
timestamp 1644511149
transform 1 0 22540 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_245
timestamp 1644511149
transform 1 0 23644 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_251
timestamp 1644511149
transform 1 0 24196 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_253
timestamp 1644511149
transform 1 0 24380 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_265
timestamp 1644511149
transform 1 0 25484 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_277
timestamp 1644511149
transform 1 0 26588 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_289
timestamp 1644511149
transform 1 0 27692 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_301
timestamp 1644511149
transform 1 0 28796 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_307
timestamp 1644511149
transform 1 0 29348 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_309
timestamp 1644511149
transform 1 0 29532 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_321
timestamp 1644511149
transform 1 0 30636 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_333
timestamp 1644511149
transform 1 0 31740 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_345
timestamp 1644511149
transform 1 0 32844 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_357
timestamp 1644511149
transform 1 0 33948 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_363
timestamp 1644511149
transform 1 0 34500 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_365
timestamp 1644511149
transform 1 0 34684 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_377
timestamp 1644511149
transform 1 0 35788 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_389
timestamp 1644511149
transform 1 0 36892 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_401
timestamp 1644511149
transform 1 0 37996 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_413
timestamp 1644511149
transform 1 0 39100 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_419
timestamp 1644511149
transform 1 0 39652 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_421
timestamp 1644511149
transform 1 0 39836 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_433
timestamp 1644511149
transform 1 0 40940 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_445
timestamp 1644511149
transform 1 0 42044 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_457
timestamp 1644511149
transform 1 0 43148 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_469
timestamp 1644511149
transform 1 0 44252 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_475
timestamp 1644511149
transform 1 0 44804 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_477
timestamp 1644511149
transform 1 0 44988 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_489
timestamp 1644511149
transform 1 0 46092 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_501
timestamp 1644511149
transform 1 0 47196 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_513
timestamp 1644511149
transform 1 0 48300 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_525
timestamp 1644511149
transform 1 0 49404 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_531
timestamp 1644511149
transform 1 0 49956 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_533
timestamp 1644511149
transform 1 0 50140 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_545
timestamp 1644511149
transform 1 0 51244 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_557
timestamp 1644511149
transform 1 0 52348 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_569
timestamp 1644511149
transform 1 0 53452 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_581
timestamp 1644511149
transform 1 0 54556 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_587
timestamp 1644511149
transform 1 0 55108 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_589
timestamp 1644511149
transform 1 0 55292 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_54_601
timestamp 1644511149
transform 1 0 56396 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_621
timestamp 1644511149
transform 1 0 58236 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_55_3
timestamp 1644511149
transform 1 0 1380 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_15
timestamp 1644511149
transform 1 0 2484 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_27
timestamp 1644511149
transform 1 0 3588 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_39
timestamp 1644511149
transform 1 0 4692 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_51
timestamp 1644511149
transform 1 0 5796 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_55
timestamp 1644511149
transform 1 0 6164 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_57
timestamp 1644511149
transform 1 0 6348 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_69
timestamp 1644511149
transform 1 0 7452 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_81
timestamp 1644511149
transform 1 0 8556 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_93
timestamp 1644511149
transform 1 0 9660 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_105
timestamp 1644511149
transform 1 0 10764 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_111
timestamp 1644511149
transform 1 0 11316 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_113
timestamp 1644511149
transform 1 0 11500 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_125
timestamp 1644511149
transform 1 0 12604 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_137
timestamp 1644511149
transform 1 0 13708 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_149
timestamp 1644511149
transform 1 0 14812 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_161
timestamp 1644511149
transform 1 0 15916 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_167
timestamp 1644511149
transform 1 0 16468 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_169
timestamp 1644511149
transform 1 0 16652 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_181
timestamp 1644511149
transform 1 0 17756 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_193
timestamp 1644511149
transform 1 0 18860 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_205
timestamp 1644511149
transform 1 0 19964 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_217
timestamp 1644511149
transform 1 0 21068 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_223
timestamp 1644511149
transform 1 0 21620 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_225
timestamp 1644511149
transform 1 0 21804 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_237
timestamp 1644511149
transform 1 0 22908 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_249
timestamp 1644511149
transform 1 0 24012 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_261
timestamp 1644511149
transform 1 0 25116 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_273
timestamp 1644511149
transform 1 0 26220 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_279
timestamp 1644511149
transform 1 0 26772 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_281
timestamp 1644511149
transform 1 0 26956 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_293
timestamp 1644511149
transform 1 0 28060 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_305
timestamp 1644511149
transform 1 0 29164 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_317
timestamp 1644511149
transform 1 0 30268 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_329
timestamp 1644511149
transform 1 0 31372 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_335
timestamp 1644511149
transform 1 0 31924 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_337
timestamp 1644511149
transform 1 0 32108 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_349
timestamp 1644511149
transform 1 0 33212 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_361
timestamp 1644511149
transform 1 0 34316 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_373
timestamp 1644511149
transform 1 0 35420 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_385
timestamp 1644511149
transform 1 0 36524 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_391
timestamp 1644511149
transform 1 0 37076 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_393
timestamp 1644511149
transform 1 0 37260 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_405
timestamp 1644511149
transform 1 0 38364 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_417
timestamp 1644511149
transform 1 0 39468 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_429
timestamp 1644511149
transform 1 0 40572 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_441
timestamp 1644511149
transform 1 0 41676 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_447
timestamp 1644511149
transform 1 0 42228 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_449
timestamp 1644511149
transform 1 0 42412 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_461
timestamp 1644511149
transform 1 0 43516 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_473
timestamp 1644511149
transform 1 0 44620 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_485
timestamp 1644511149
transform 1 0 45724 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_497
timestamp 1644511149
transform 1 0 46828 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_503
timestamp 1644511149
transform 1 0 47380 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_505
timestamp 1644511149
transform 1 0 47564 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_517
timestamp 1644511149
transform 1 0 48668 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_529
timestamp 1644511149
transform 1 0 49772 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_541
timestamp 1644511149
transform 1 0 50876 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_553
timestamp 1644511149
transform 1 0 51980 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_559
timestamp 1644511149
transform 1 0 52532 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_561
timestamp 1644511149
transform 1 0 52716 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_573
timestamp 1644511149
transform 1 0 53820 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_585
timestamp 1644511149
transform 1 0 54924 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_597
timestamp 1644511149
transform 1 0 56028 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_609
timestamp 1644511149
transform 1 0 57132 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_615
timestamp 1644511149
transform 1 0 57684 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_55_617
timestamp 1644511149
transform 1 0 57868 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_56_3
timestamp 1644511149
transform 1 0 1380 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_15
timestamp 1644511149
transform 1 0 2484 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_56_27
timestamp 1644511149
transform 1 0 3588 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_29
timestamp 1644511149
transform 1 0 3772 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_41
timestamp 1644511149
transform 1 0 4876 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_53
timestamp 1644511149
transform 1 0 5980 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_65
timestamp 1644511149
transform 1 0 7084 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_77
timestamp 1644511149
transform 1 0 8188 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_83
timestamp 1644511149
transform 1 0 8740 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_85
timestamp 1644511149
transform 1 0 8924 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_97
timestamp 1644511149
transform 1 0 10028 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_109
timestamp 1644511149
transform 1 0 11132 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_121
timestamp 1644511149
transform 1 0 12236 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_133
timestamp 1644511149
transform 1 0 13340 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_139
timestamp 1644511149
transform 1 0 13892 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_141
timestamp 1644511149
transform 1 0 14076 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_153
timestamp 1644511149
transform 1 0 15180 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_165
timestamp 1644511149
transform 1 0 16284 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_177
timestamp 1644511149
transform 1 0 17388 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_189
timestamp 1644511149
transform 1 0 18492 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_195
timestamp 1644511149
transform 1 0 19044 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_197
timestamp 1644511149
transform 1 0 19228 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_209
timestamp 1644511149
transform 1 0 20332 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_221
timestamp 1644511149
transform 1 0 21436 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_233
timestamp 1644511149
transform 1 0 22540 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_245
timestamp 1644511149
transform 1 0 23644 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_251
timestamp 1644511149
transform 1 0 24196 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_253
timestamp 1644511149
transform 1 0 24380 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_265
timestamp 1644511149
transform 1 0 25484 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_277
timestamp 1644511149
transform 1 0 26588 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_289
timestamp 1644511149
transform 1 0 27692 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_301
timestamp 1644511149
transform 1 0 28796 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_307
timestamp 1644511149
transform 1 0 29348 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_309
timestamp 1644511149
transform 1 0 29532 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_321
timestamp 1644511149
transform 1 0 30636 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_333
timestamp 1644511149
transform 1 0 31740 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_345
timestamp 1644511149
transform 1 0 32844 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_357
timestamp 1644511149
transform 1 0 33948 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_363
timestamp 1644511149
transform 1 0 34500 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_365
timestamp 1644511149
transform 1 0 34684 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_377
timestamp 1644511149
transform 1 0 35788 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_389
timestamp 1644511149
transform 1 0 36892 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_401
timestamp 1644511149
transform 1 0 37996 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_413
timestamp 1644511149
transform 1 0 39100 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_419
timestamp 1644511149
transform 1 0 39652 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_421
timestamp 1644511149
transform 1 0 39836 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_433
timestamp 1644511149
transform 1 0 40940 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_445
timestamp 1644511149
transform 1 0 42044 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_457
timestamp 1644511149
transform 1 0 43148 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_469
timestamp 1644511149
transform 1 0 44252 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_475
timestamp 1644511149
transform 1 0 44804 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_477
timestamp 1644511149
transform 1 0 44988 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_489
timestamp 1644511149
transform 1 0 46092 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_501
timestamp 1644511149
transform 1 0 47196 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_513
timestamp 1644511149
transform 1 0 48300 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_525
timestamp 1644511149
transform 1 0 49404 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_531
timestamp 1644511149
transform 1 0 49956 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_533
timestamp 1644511149
transform 1 0 50140 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_545
timestamp 1644511149
transform 1 0 51244 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_557
timestamp 1644511149
transform 1 0 52348 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_569
timestamp 1644511149
transform 1 0 53452 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_581
timestamp 1644511149
transform 1 0 54556 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_587
timestamp 1644511149
transform 1 0 55108 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_589
timestamp 1644511149
transform 1 0 55292 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_601
timestamp 1644511149
transform 1 0 56396 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_613
timestamp 1644511149
transform 1 0 57500 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_3
timestamp 1644511149
transform 1 0 1380 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_15
timestamp 1644511149
transform 1 0 2484 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_27
timestamp 1644511149
transform 1 0 3588 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_39
timestamp 1644511149
transform 1 0 4692 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_51
timestamp 1644511149
transform 1 0 5796 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_55
timestamp 1644511149
transform 1 0 6164 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_57
timestamp 1644511149
transform 1 0 6348 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_69
timestamp 1644511149
transform 1 0 7452 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_81
timestamp 1644511149
transform 1 0 8556 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_93
timestamp 1644511149
transform 1 0 9660 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_105
timestamp 1644511149
transform 1 0 10764 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_111
timestamp 1644511149
transform 1 0 11316 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_113
timestamp 1644511149
transform 1 0 11500 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_125
timestamp 1644511149
transform 1 0 12604 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_137
timestamp 1644511149
transform 1 0 13708 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_149
timestamp 1644511149
transform 1 0 14812 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_161
timestamp 1644511149
transform 1 0 15916 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_167
timestamp 1644511149
transform 1 0 16468 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_169
timestamp 1644511149
transform 1 0 16652 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_181
timestamp 1644511149
transform 1 0 17756 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_193
timestamp 1644511149
transform 1 0 18860 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_205
timestamp 1644511149
transform 1 0 19964 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_217
timestamp 1644511149
transform 1 0 21068 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_223
timestamp 1644511149
transform 1 0 21620 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_225
timestamp 1644511149
transform 1 0 21804 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_237
timestamp 1644511149
transform 1 0 22908 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_249
timestamp 1644511149
transform 1 0 24012 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_261
timestamp 1644511149
transform 1 0 25116 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_273
timestamp 1644511149
transform 1 0 26220 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_279
timestamp 1644511149
transform 1 0 26772 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_281
timestamp 1644511149
transform 1 0 26956 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_293
timestamp 1644511149
transform 1 0 28060 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_305
timestamp 1644511149
transform 1 0 29164 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_317
timestamp 1644511149
transform 1 0 30268 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_329
timestamp 1644511149
transform 1 0 31372 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_335
timestamp 1644511149
transform 1 0 31924 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_337
timestamp 1644511149
transform 1 0 32108 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_349
timestamp 1644511149
transform 1 0 33212 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_361
timestamp 1644511149
transform 1 0 34316 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_373
timestamp 1644511149
transform 1 0 35420 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_385
timestamp 1644511149
transform 1 0 36524 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_391
timestamp 1644511149
transform 1 0 37076 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_393
timestamp 1644511149
transform 1 0 37260 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_405
timestamp 1644511149
transform 1 0 38364 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_417
timestamp 1644511149
transform 1 0 39468 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_429
timestamp 1644511149
transform 1 0 40572 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_441
timestamp 1644511149
transform 1 0 41676 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_447
timestamp 1644511149
transform 1 0 42228 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_449
timestamp 1644511149
transform 1 0 42412 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_461
timestamp 1644511149
transform 1 0 43516 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_473
timestamp 1644511149
transform 1 0 44620 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_485
timestamp 1644511149
transform 1 0 45724 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_497
timestamp 1644511149
transform 1 0 46828 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_503
timestamp 1644511149
transform 1 0 47380 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_505
timestamp 1644511149
transform 1 0 47564 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_517
timestamp 1644511149
transform 1 0 48668 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_529
timestamp 1644511149
transform 1 0 49772 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_541
timestamp 1644511149
transform 1 0 50876 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_553
timestamp 1644511149
transform 1 0 51980 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_559
timestamp 1644511149
transform 1 0 52532 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_561
timestamp 1644511149
transform 1 0 52716 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_573
timestamp 1644511149
transform 1 0 53820 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_585
timestamp 1644511149
transform 1 0 54924 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_597
timestamp 1644511149
transform 1 0 56028 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_609
timestamp 1644511149
transform 1 0 57132 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_615
timestamp 1644511149
transform 1 0 57684 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_57_617
timestamp 1644511149
transform 1 0 57868 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_58_3
timestamp 1644511149
transform 1 0 1380 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_15
timestamp 1644511149
transform 1 0 2484 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_58_27
timestamp 1644511149
transform 1 0 3588 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_29
timestamp 1644511149
transform 1 0 3772 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_41
timestamp 1644511149
transform 1 0 4876 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_53
timestamp 1644511149
transform 1 0 5980 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_65
timestamp 1644511149
transform 1 0 7084 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_77
timestamp 1644511149
transform 1 0 8188 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_83
timestamp 1644511149
transform 1 0 8740 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_85
timestamp 1644511149
transform 1 0 8924 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_97
timestamp 1644511149
transform 1 0 10028 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_109
timestamp 1644511149
transform 1 0 11132 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_121
timestamp 1644511149
transform 1 0 12236 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_133
timestamp 1644511149
transform 1 0 13340 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_139
timestamp 1644511149
transform 1 0 13892 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_141
timestamp 1644511149
transform 1 0 14076 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_153
timestamp 1644511149
transform 1 0 15180 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_165
timestamp 1644511149
transform 1 0 16284 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_177
timestamp 1644511149
transform 1 0 17388 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_189
timestamp 1644511149
transform 1 0 18492 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_195
timestamp 1644511149
transform 1 0 19044 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_197
timestamp 1644511149
transform 1 0 19228 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_209
timestamp 1644511149
transform 1 0 20332 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_221
timestamp 1644511149
transform 1 0 21436 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_233
timestamp 1644511149
transform 1 0 22540 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_245
timestamp 1644511149
transform 1 0 23644 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_251
timestamp 1644511149
transform 1 0 24196 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_253
timestamp 1644511149
transform 1 0 24380 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_265
timestamp 1644511149
transform 1 0 25484 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_277
timestamp 1644511149
transform 1 0 26588 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_289
timestamp 1644511149
transform 1 0 27692 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_301
timestamp 1644511149
transform 1 0 28796 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_307
timestamp 1644511149
transform 1 0 29348 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_309
timestamp 1644511149
transform 1 0 29532 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_321
timestamp 1644511149
transform 1 0 30636 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_333
timestamp 1644511149
transform 1 0 31740 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_345
timestamp 1644511149
transform 1 0 32844 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_357
timestamp 1644511149
transform 1 0 33948 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_363
timestamp 1644511149
transform 1 0 34500 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_365
timestamp 1644511149
transform 1 0 34684 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_377
timestamp 1644511149
transform 1 0 35788 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_389
timestamp 1644511149
transform 1 0 36892 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_401
timestamp 1644511149
transform 1 0 37996 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_413
timestamp 1644511149
transform 1 0 39100 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_419
timestamp 1644511149
transform 1 0 39652 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_421
timestamp 1644511149
transform 1 0 39836 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_433
timestamp 1644511149
transform 1 0 40940 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_445
timestamp 1644511149
transform 1 0 42044 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_457
timestamp 1644511149
transform 1 0 43148 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_469
timestamp 1644511149
transform 1 0 44252 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_475
timestamp 1644511149
transform 1 0 44804 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_477
timestamp 1644511149
transform 1 0 44988 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_489
timestamp 1644511149
transform 1 0 46092 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_501
timestamp 1644511149
transform 1 0 47196 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_513
timestamp 1644511149
transform 1 0 48300 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_525
timestamp 1644511149
transform 1 0 49404 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_531
timestamp 1644511149
transform 1 0 49956 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_533
timestamp 1644511149
transform 1 0 50140 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_545
timestamp 1644511149
transform 1 0 51244 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_557
timestamp 1644511149
transform 1 0 52348 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_569
timestamp 1644511149
transform 1 0 53452 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_581
timestamp 1644511149
transform 1 0 54556 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_587
timestamp 1644511149
transform 1 0 55108 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_589
timestamp 1644511149
transform 1 0 55292 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_601
timestamp 1644511149
transform 1 0 56396 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_613
timestamp 1644511149
transform 1 0 57500 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_59_3
timestamp 1644511149
transform 1 0 1380 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_59_32
timestamp 1644511149
transform 1 0 4048 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_44
timestamp 1644511149
transform 1 0 5152 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_57
timestamp 1644511149
transform 1 0 6348 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_69
timestamp 1644511149
transform 1 0 7452 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_81
timestamp 1644511149
transform 1 0 8556 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_93
timestamp 1644511149
transform 1 0 9660 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_105
timestamp 1644511149
transform 1 0 10764 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_111
timestamp 1644511149
transform 1 0 11316 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_113
timestamp 1644511149
transform 1 0 11500 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_125
timestamp 1644511149
transform 1 0 12604 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_137
timestamp 1644511149
transform 1 0 13708 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_149
timestamp 1644511149
transform 1 0 14812 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_161
timestamp 1644511149
transform 1 0 15916 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_167
timestamp 1644511149
transform 1 0 16468 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_169
timestamp 1644511149
transform 1 0 16652 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_181
timestamp 1644511149
transform 1 0 17756 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_193
timestamp 1644511149
transform 1 0 18860 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_205
timestamp 1644511149
transform 1 0 19964 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_217
timestamp 1644511149
transform 1 0 21068 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_223
timestamp 1644511149
transform 1 0 21620 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_225
timestamp 1644511149
transform 1 0 21804 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_237
timestamp 1644511149
transform 1 0 22908 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_249
timestamp 1644511149
transform 1 0 24012 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_261
timestamp 1644511149
transform 1 0 25116 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_273
timestamp 1644511149
transform 1 0 26220 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_279
timestamp 1644511149
transform 1 0 26772 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_281
timestamp 1644511149
transform 1 0 26956 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_293
timestamp 1644511149
transform 1 0 28060 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_305
timestamp 1644511149
transform 1 0 29164 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_317
timestamp 1644511149
transform 1 0 30268 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_329
timestamp 1644511149
transform 1 0 31372 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_335
timestamp 1644511149
transform 1 0 31924 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_337
timestamp 1644511149
transform 1 0 32108 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_349
timestamp 1644511149
transform 1 0 33212 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_361
timestamp 1644511149
transform 1 0 34316 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_373
timestamp 1644511149
transform 1 0 35420 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_385
timestamp 1644511149
transform 1 0 36524 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_391
timestamp 1644511149
transform 1 0 37076 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_393
timestamp 1644511149
transform 1 0 37260 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_405
timestamp 1644511149
transform 1 0 38364 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_417
timestamp 1644511149
transform 1 0 39468 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_429
timestamp 1644511149
transform 1 0 40572 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_441
timestamp 1644511149
transform 1 0 41676 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_447
timestamp 1644511149
transform 1 0 42228 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_449
timestamp 1644511149
transform 1 0 42412 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_461
timestamp 1644511149
transform 1 0 43516 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_473
timestamp 1644511149
transform 1 0 44620 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_485
timestamp 1644511149
transform 1 0 45724 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_497
timestamp 1644511149
transform 1 0 46828 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_503
timestamp 1644511149
transform 1 0 47380 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_505
timestamp 1644511149
transform 1 0 47564 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_517
timestamp 1644511149
transform 1 0 48668 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_529
timestamp 1644511149
transform 1 0 49772 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_541
timestamp 1644511149
transform 1 0 50876 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_553
timestamp 1644511149
transform 1 0 51980 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_559
timestamp 1644511149
transform 1 0 52532 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_561
timestamp 1644511149
transform 1 0 52716 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_573
timestamp 1644511149
transform 1 0 53820 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_585
timestamp 1644511149
transform 1 0 54924 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_597
timestamp 1644511149
transform 1 0 56028 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_609
timestamp 1644511149
transform 1 0 57132 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_615
timestamp 1644511149
transform 1 0 57684 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_59_617
timestamp 1644511149
transform 1 0 57868 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_60_3
timestamp 1644511149
transform 1 0 1380 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_60_11
timestamp 1644511149
transform 1 0 2116 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_15
timestamp 1644511149
transform 1 0 2484 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_60_27
timestamp 1644511149
transform 1 0 3588 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_32
timestamp 1644511149
transform 1 0 4048 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_44
timestamp 1644511149
transform 1 0 5152 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_56
timestamp 1644511149
transform 1 0 6256 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_68
timestamp 1644511149
transform 1 0 7360 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_60_80
timestamp 1644511149
transform 1 0 8464 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_60_85
timestamp 1644511149
transform 1 0 8924 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_97
timestamp 1644511149
transform 1 0 10028 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_109
timestamp 1644511149
transform 1 0 11132 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_121
timestamp 1644511149
transform 1 0 12236 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_133
timestamp 1644511149
transform 1 0 13340 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_139
timestamp 1644511149
transform 1 0 13892 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_141
timestamp 1644511149
transform 1 0 14076 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_153
timestamp 1644511149
transform 1 0 15180 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_165
timestamp 1644511149
transform 1 0 16284 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_177
timestamp 1644511149
transform 1 0 17388 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_189
timestamp 1644511149
transform 1 0 18492 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_195
timestamp 1644511149
transform 1 0 19044 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_197
timestamp 1644511149
transform 1 0 19228 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_209
timestamp 1644511149
transform 1 0 20332 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_221
timestamp 1644511149
transform 1 0 21436 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_233
timestamp 1644511149
transform 1 0 22540 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_245
timestamp 1644511149
transform 1 0 23644 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_251
timestamp 1644511149
transform 1 0 24196 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_253
timestamp 1644511149
transform 1 0 24380 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_265
timestamp 1644511149
transform 1 0 25484 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_277
timestamp 1644511149
transform 1 0 26588 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_289
timestamp 1644511149
transform 1 0 27692 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_301
timestamp 1644511149
transform 1 0 28796 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_307
timestamp 1644511149
transform 1 0 29348 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_309
timestamp 1644511149
transform 1 0 29532 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_321
timestamp 1644511149
transform 1 0 30636 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_333
timestamp 1644511149
transform 1 0 31740 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_345
timestamp 1644511149
transform 1 0 32844 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_357
timestamp 1644511149
transform 1 0 33948 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_363
timestamp 1644511149
transform 1 0 34500 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_365
timestamp 1644511149
transform 1 0 34684 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_377
timestamp 1644511149
transform 1 0 35788 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_389
timestamp 1644511149
transform 1 0 36892 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_401
timestamp 1644511149
transform 1 0 37996 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_413
timestamp 1644511149
transform 1 0 39100 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_419
timestamp 1644511149
transform 1 0 39652 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_421
timestamp 1644511149
transform 1 0 39836 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_433
timestamp 1644511149
transform 1 0 40940 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_445
timestamp 1644511149
transform 1 0 42044 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_457
timestamp 1644511149
transform 1 0 43148 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_469
timestamp 1644511149
transform 1 0 44252 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_475
timestamp 1644511149
transform 1 0 44804 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_477
timestamp 1644511149
transform 1 0 44988 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_489
timestamp 1644511149
transform 1 0 46092 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_501
timestamp 1644511149
transform 1 0 47196 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_513
timestamp 1644511149
transform 1 0 48300 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_525
timestamp 1644511149
transform 1 0 49404 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_531
timestamp 1644511149
transform 1 0 49956 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_533
timestamp 1644511149
transform 1 0 50140 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_545
timestamp 1644511149
transform 1 0 51244 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_557
timestamp 1644511149
transform 1 0 52348 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_569
timestamp 1644511149
transform 1 0 53452 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_581
timestamp 1644511149
transform 1 0 54556 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_587
timestamp 1644511149
transform 1 0 55108 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_589
timestamp 1644511149
transform 1 0 55292 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_601
timestamp 1644511149
transform 1 0 56396 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_613
timestamp 1644511149
transform 1 0 57500 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_3
timestamp 1644511149
transform 1 0 1380 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_15
timestamp 1644511149
transform 1 0 2484 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_27
timestamp 1644511149
transform 1 0 3588 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_39
timestamp 1644511149
transform 1 0 4692 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_61_51
timestamp 1644511149
transform 1 0 5796 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_55
timestamp 1644511149
transform 1 0 6164 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_57
timestamp 1644511149
transform 1 0 6348 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_69
timestamp 1644511149
transform 1 0 7452 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_81
timestamp 1644511149
transform 1 0 8556 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_93
timestamp 1644511149
transform 1 0 9660 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_105
timestamp 1644511149
transform 1 0 10764 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_111
timestamp 1644511149
transform 1 0 11316 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_113
timestamp 1644511149
transform 1 0 11500 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_125
timestamp 1644511149
transform 1 0 12604 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_137
timestamp 1644511149
transform 1 0 13708 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_149
timestamp 1644511149
transform 1 0 14812 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_161
timestamp 1644511149
transform 1 0 15916 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_167
timestamp 1644511149
transform 1 0 16468 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_169
timestamp 1644511149
transform 1 0 16652 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_181
timestamp 1644511149
transform 1 0 17756 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_193
timestamp 1644511149
transform 1 0 18860 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_205
timestamp 1644511149
transform 1 0 19964 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_217
timestamp 1644511149
transform 1 0 21068 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_223
timestamp 1644511149
transform 1 0 21620 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_225
timestamp 1644511149
transform 1 0 21804 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_237
timestamp 1644511149
transform 1 0 22908 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_249
timestamp 1644511149
transform 1 0 24012 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_261
timestamp 1644511149
transform 1 0 25116 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_273
timestamp 1644511149
transform 1 0 26220 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_279
timestamp 1644511149
transform 1 0 26772 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_281
timestamp 1644511149
transform 1 0 26956 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_293
timestamp 1644511149
transform 1 0 28060 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_305
timestamp 1644511149
transform 1 0 29164 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_317
timestamp 1644511149
transform 1 0 30268 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_329
timestamp 1644511149
transform 1 0 31372 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_335
timestamp 1644511149
transform 1 0 31924 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_337
timestamp 1644511149
transform 1 0 32108 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_349
timestamp 1644511149
transform 1 0 33212 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_361
timestamp 1644511149
transform 1 0 34316 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_373
timestamp 1644511149
transform 1 0 35420 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_385
timestamp 1644511149
transform 1 0 36524 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_391
timestamp 1644511149
transform 1 0 37076 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_393
timestamp 1644511149
transform 1 0 37260 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_405
timestamp 1644511149
transform 1 0 38364 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_417
timestamp 1644511149
transform 1 0 39468 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_429
timestamp 1644511149
transform 1 0 40572 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_441
timestamp 1644511149
transform 1 0 41676 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_447
timestamp 1644511149
transform 1 0 42228 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_449
timestamp 1644511149
transform 1 0 42412 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_461
timestamp 1644511149
transform 1 0 43516 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_473
timestamp 1644511149
transform 1 0 44620 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_485
timestamp 1644511149
transform 1 0 45724 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_497
timestamp 1644511149
transform 1 0 46828 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_503
timestamp 1644511149
transform 1 0 47380 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_505
timestamp 1644511149
transform 1 0 47564 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_517
timestamp 1644511149
transform 1 0 48668 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_529
timestamp 1644511149
transform 1 0 49772 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_541
timestamp 1644511149
transform 1 0 50876 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_553
timestamp 1644511149
transform 1 0 51980 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_559
timestamp 1644511149
transform 1 0 52532 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_561
timestamp 1644511149
transform 1 0 52716 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_573
timestamp 1644511149
transform 1 0 53820 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_585
timestamp 1644511149
transform 1 0 54924 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_597
timestamp 1644511149
transform 1 0 56028 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_609
timestamp 1644511149
transform 1 0 57132 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_615
timestamp 1644511149
transform 1 0 57684 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_61_617
timestamp 1644511149
transform 1 0 57868 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_62_3
timestamp 1644511149
transform 1 0 1380 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_15
timestamp 1644511149
transform 1 0 2484 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_62_27
timestamp 1644511149
transform 1 0 3588 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_29
timestamp 1644511149
transform 1 0 3772 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_41
timestamp 1644511149
transform 1 0 4876 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_53
timestamp 1644511149
transform 1 0 5980 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_65
timestamp 1644511149
transform 1 0 7084 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_77
timestamp 1644511149
transform 1 0 8188 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_83
timestamp 1644511149
transform 1 0 8740 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_85
timestamp 1644511149
transform 1 0 8924 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_97
timestamp 1644511149
transform 1 0 10028 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_109
timestamp 1644511149
transform 1 0 11132 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_121
timestamp 1644511149
transform 1 0 12236 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_133
timestamp 1644511149
transform 1 0 13340 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_139
timestamp 1644511149
transform 1 0 13892 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_141
timestamp 1644511149
transform 1 0 14076 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_153
timestamp 1644511149
transform 1 0 15180 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_165
timestamp 1644511149
transform 1 0 16284 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_177
timestamp 1644511149
transform 1 0 17388 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_189
timestamp 1644511149
transform 1 0 18492 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_195
timestamp 1644511149
transform 1 0 19044 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_197
timestamp 1644511149
transform 1 0 19228 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_209
timestamp 1644511149
transform 1 0 20332 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_221
timestamp 1644511149
transform 1 0 21436 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_233
timestamp 1644511149
transform 1 0 22540 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_245
timestamp 1644511149
transform 1 0 23644 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_251
timestamp 1644511149
transform 1 0 24196 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_253
timestamp 1644511149
transform 1 0 24380 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_265
timestamp 1644511149
transform 1 0 25484 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_277
timestamp 1644511149
transform 1 0 26588 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_289
timestamp 1644511149
transform 1 0 27692 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_301
timestamp 1644511149
transform 1 0 28796 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_307
timestamp 1644511149
transform 1 0 29348 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_309
timestamp 1644511149
transform 1 0 29532 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_321
timestamp 1644511149
transform 1 0 30636 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_333
timestamp 1644511149
transform 1 0 31740 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_345
timestamp 1644511149
transform 1 0 32844 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_357
timestamp 1644511149
transform 1 0 33948 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_363
timestamp 1644511149
transform 1 0 34500 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_365
timestamp 1644511149
transform 1 0 34684 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_377
timestamp 1644511149
transform 1 0 35788 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_389
timestamp 1644511149
transform 1 0 36892 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_401
timestamp 1644511149
transform 1 0 37996 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_413
timestamp 1644511149
transform 1 0 39100 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_419
timestamp 1644511149
transform 1 0 39652 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_421
timestamp 1644511149
transform 1 0 39836 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_433
timestamp 1644511149
transform 1 0 40940 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_445
timestamp 1644511149
transform 1 0 42044 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_457
timestamp 1644511149
transform 1 0 43148 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_469
timestamp 1644511149
transform 1 0 44252 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_475
timestamp 1644511149
transform 1 0 44804 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_477
timestamp 1644511149
transform 1 0 44988 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_489
timestamp 1644511149
transform 1 0 46092 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_501
timestamp 1644511149
transform 1 0 47196 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_513
timestamp 1644511149
transform 1 0 48300 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_525
timestamp 1644511149
transform 1 0 49404 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_531
timestamp 1644511149
transform 1 0 49956 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_533
timestamp 1644511149
transform 1 0 50140 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_545
timestamp 1644511149
transform 1 0 51244 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_557
timestamp 1644511149
transform 1 0 52348 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_569
timestamp 1644511149
transform 1 0 53452 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_581
timestamp 1644511149
transform 1 0 54556 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_587
timestamp 1644511149
transform 1 0 55108 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_589
timestamp 1644511149
transform 1 0 55292 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_601
timestamp 1644511149
transform 1 0 56396 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_613
timestamp 1644511149
transform 1 0 57500 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_3
timestamp 1644511149
transform 1 0 1380 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_15
timestamp 1644511149
transform 1 0 2484 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_27
timestamp 1644511149
transform 1 0 3588 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_39
timestamp 1644511149
transform 1 0 4692 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_63_51
timestamp 1644511149
transform 1 0 5796 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_55
timestamp 1644511149
transform 1 0 6164 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_57
timestamp 1644511149
transform 1 0 6348 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_69
timestamp 1644511149
transform 1 0 7452 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_81
timestamp 1644511149
transform 1 0 8556 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_93
timestamp 1644511149
transform 1 0 9660 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_105
timestamp 1644511149
transform 1 0 10764 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_111
timestamp 1644511149
transform 1 0 11316 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_113
timestamp 1644511149
transform 1 0 11500 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_125
timestamp 1644511149
transform 1 0 12604 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_137
timestamp 1644511149
transform 1 0 13708 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_149
timestamp 1644511149
transform 1 0 14812 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_161
timestamp 1644511149
transform 1 0 15916 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_167
timestamp 1644511149
transform 1 0 16468 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_169
timestamp 1644511149
transform 1 0 16652 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_181
timestamp 1644511149
transform 1 0 17756 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_193
timestamp 1644511149
transform 1 0 18860 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_205
timestamp 1644511149
transform 1 0 19964 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_217
timestamp 1644511149
transform 1 0 21068 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_223
timestamp 1644511149
transform 1 0 21620 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_225
timestamp 1644511149
transform 1 0 21804 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_237
timestamp 1644511149
transform 1 0 22908 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_249
timestamp 1644511149
transform 1 0 24012 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_261
timestamp 1644511149
transform 1 0 25116 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_273
timestamp 1644511149
transform 1 0 26220 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_279
timestamp 1644511149
transform 1 0 26772 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_281
timestamp 1644511149
transform 1 0 26956 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_293
timestamp 1644511149
transform 1 0 28060 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_305
timestamp 1644511149
transform 1 0 29164 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_317
timestamp 1644511149
transform 1 0 30268 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_329
timestamp 1644511149
transform 1 0 31372 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_335
timestamp 1644511149
transform 1 0 31924 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_337
timestamp 1644511149
transform 1 0 32108 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_349
timestamp 1644511149
transform 1 0 33212 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_361
timestamp 1644511149
transform 1 0 34316 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_373
timestamp 1644511149
transform 1 0 35420 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_385
timestamp 1644511149
transform 1 0 36524 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_391
timestamp 1644511149
transform 1 0 37076 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_393
timestamp 1644511149
transform 1 0 37260 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_405
timestamp 1644511149
transform 1 0 38364 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_417
timestamp 1644511149
transform 1 0 39468 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_429
timestamp 1644511149
transform 1 0 40572 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_441
timestamp 1644511149
transform 1 0 41676 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_447
timestamp 1644511149
transform 1 0 42228 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_449
timestamp 1644511149
transform 1 0 42412 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_461
timestamp 1644511149
transform 1 0 43516 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_473
timestamp 1644511149
transform 1 0 44620 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_485
timestamp 1644511149
transform 1 0 45724 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_497
timestamp 1644511149
transform 1 0 46828 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_503
timestamp 1644511149
transform 1 0 47380 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_505
timestamp 1644511149
transform 1 0 47564 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_517
timestamp 1644511149
transform 1 0 48668 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_529
timestamp 1644511149
transform 1 0 49772 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_541
timestamp 1644511149
transform 1 0 50876 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_553
timestamp 1644511149
transform 1 0 51980 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_559
timestamp 1644511149
transform 1 0 52532 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_561
timestamp 1644511149
transform 1 0 52716 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_573
timestamp 1644511149
transform 1 0 53820 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_585
timestamp 1644511149
transform 1 0 54924 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_597
timestamp 1644511149
transform 1 0 56028 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_609
timestamp 1644511149
transform 1 0 57132 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_615
timestamp 1644511149
transform 1 0 57684 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_63_617
timestamp 1644511149
transform 1 0 57868 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_64_3
timestamp 1644511149
transform 1 0 1380 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_15
timestamp 1644511149
transform 1 0 2484 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_64_27
timestamp 1644511149
transform 1 0 3588 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_29
timestamp 1644511149
transform 1 0 3772 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_41
timestamp 1644511149
transform 1 0 4876 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_53
timestamp 1644511149
transform 1 0 5980 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_65
timestamp 1644511149
transform 1 0 7084 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_77
timestamp 1644511149
transform 1 0 8188 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_83
timestamp 1644511149
transform 1 0 8740 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_85
timestamp 1644511149
transform 1 0 8924 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_97
timestamp 1644511149
transform 1 0 10028 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_109
timestamp 1644511149
transform 1 0 11132 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_121
timestamp 1644511149
transform 1 0 12236 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_133
timestamp 1644511149
transform 1 0 13340 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_139
timestamp 1644511149
transform 1 0 13892 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_141
timestamp 1644511149
transform 1 0 14076 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_153
timestamp 1644511149
transform 1 0 15180 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_165
timestamp 1644511149
transform 1 0 16284 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_177
timestamp 1644511149
transform 1 0 17388 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_189
timestamp 1644511149
transform 1 0 18492 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_195
timestamp 1644511149
transform 1 0 19044 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_197
timestamp 1644511149
transform 1 0 19228 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_209
timestamp 1644511149
transform 1 0 20332 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_221
timestamp 1644511149
transform 1 0 21436 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_233
timestamp 1644511149
transform 1 0 22540 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_245
timestamp 1644511149
transform 1 0 23644 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_251
timestamp 1644511149
transform 1 0 24196 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_253
timestamp 1644511149
transform 1 0 24380 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_265
timestamp 1644511149
transform 1 0 25484 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_277
timestamp 1644511149
transform 1 0 26588 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_289
timestamp 1644511149
transform 1 0 27692 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_301
timestamp 1644511149
transform 1 0 28796 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_307
timestamp 1644511149
transform 1 0 29348 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_309
timestamp 1644511149
transform 1 0 29532 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_321
timestamp 1644511149
transform 1 0 30636 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_333
timestamp 1644511149
transform 1 0 31740 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_345
timestamp 1644511149
transform 1 0 32844 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_357
timestamp 1644511149
transform 1 0 33948 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_363
timestamp 1644511149
transform 1 0 34500 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_365
timestamp 1644511149
transform 1 0 34684 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_377
timestamp 1644511149
transform 1 0 35788 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_389
timestamp 1644511149
transform 1 0 36892 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_401
timestamp 1644511149
transform 1 0 37996 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_413
timestamp 1644511149
transform 1 0 39100 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_419
timestamp 1644511149
transform 1 0 39652 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_421
timestamp 1644511149
transform 1 0 39836 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_433
timestamp 1644511149
transform 1 0 40940 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_445
timestamp 1644511149
transform 1 0 42044 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_457
timestamp 1644511149
transform 1 0 43148 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_469
timestamp 1644511149
transform 1 0 44252 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_475
timestamp 1644511149
transform 1 0 44804 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_477
timestamp 1644511149
transform 1 0 44988 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_489
timestamp 1644511149
transform 1 0 46092 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_501
timestamp 1644511149
transform 1 0 47196 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_513
timestamp 1644511149
transform 1 0 48300 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_525
timestamp 1644511149
transform 1 0 49404 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_531
timestamp 1644511149
transform 1 0 49956 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_533
timestamp 1644511149
transform 1 0 50140 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_545
timestamp 1644511149
transform 1 0 51244 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_557
timestamp 1644511149
transform 1 0 52348 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_569
timestamp 1644511149
transform 1 0 53452 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_581
timestamp 1644511149
transform 1 0 54556 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_587
timestamp 1644511149
transform 1 0 55108 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_589
timestamp 1644511149
transform 1 0 55292 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_601
timestamp 1644511149
transform 1 0 56396 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_613
timestamp 1644511149
transform 1 0 57500 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_3
timestamp 1644511149
transform 1 0 1380 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_15
timestamp 1644511149
transform 1 0 2484 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_27
timestamp 1644511149
transform 1 0 3588 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_39
timestamp 1644511149
transform 1 0 4692 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_65_51
timestamp 1644511149
transform 1 0 5796 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_65_55
timestamp 1644511149
transform 1 0 6164 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_57
timestamp 1644511149
transform 1 0 6348 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_69
timestamp 1644511149
transform 1 0 7452 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_81
timestamp 1644511149
transform 1 0 8556 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_93
timestamp 1644511149
transform 1 0 9660 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_105
timestamp 1644511149
transform 1 0 10764 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_111
timestamp 1644511149
transform 1 0 11316 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_113
timestamp 1644511149
transform 1 0 11500 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_125
timestamp 1644511149
transform 1 0 12604 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_137
timestamp 1644511149
transform 1 0 13708 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_149
timestamp 1644511149
transform 1 0 14812 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_161
timestamp 1644511149
transform 1 0 15916 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_167
timestamp 1644511149
transform 1 0 16468 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_169
timestamp 1644511149
transform 1 0 16652 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_181
timestamp 1644511149
transform 1 0 17756 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_193
timestamp 1644511149
transform 1 0 18860 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_205
timestamp 1644511149
transform 1 0 19964 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_217
timestamp 1644511149
transform 1 0 21068 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_223
timestamp 1644511149
transform 1 0 21620 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_225
timestamp 1644511149
transform 1 0 21804 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_237
timestamp 1644511149
transform 1 0 22908 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_249
timestamp 1644511149
transform 1 0 24012 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_261
timestamp 1644511149
transform 1 0 25116 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_273
timestamp 1644511149
transform 1 0 26220 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_279
timestamp 1644511149
transform 1 0 26772 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_281
timestamp 1644511149
transform 1 0 26956 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_293
timestamp 1644511149
transform 1 0 28060 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_305
timestamp 1644511149
transform 1 0 29164 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_317
timestamp 1644511149
transform 1 0 30268 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_329
timestamp 1644511149
transform 1 0 31372 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_335
timestamp 1644511149
transform 1 0 31924 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_337
timestamp 1644511149
transform 1 0 32108 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_349
timestamp 1644511149
transform 1 0 33212 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_361
timestamp 1644511149
transform 1 0 34316 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_373
timestamp 1644511149
transform 1 0 35420 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_385
timestamp 1644511149
transform 1 0 36524 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_391
timestamp 1644511149
transform 1 0 37076 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_393
timestamp 1644511149
transform 1 0 37260 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_405
timestamp 1644511149
transform 1 0 38364 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_417
timestamp 1644511149
transform 1 0 39468 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_429
timestamp 1644511149
transform 1 0 40572 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_441
timestamp 1644511149
transform 1 0 41676 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_447
timestamp 1644511149
transform 1 0 42228 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_449
timestamp 1644511149
transform 1 0 42412 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_461
timestamp 1644511149
transform 1 0 43516 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_473
timestamp 1644511149
transform 1 0 44620 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_485
timestamp 1644511149
transform 1 0 45724 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_497
timestamp 1644511149
transform 1 0 46828 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_503
timestamp 1644511149
transform 1 0 47380 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_505
timestamp 1644511149
transform 1 0 47564 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_517
timestamp 1644511149
transform 1 0 48668 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_529
timestamp 1644511149
transform 1 0 49772 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_541
timestamp 1644511149
transform 1 0 50876 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_553
timestamp 1644511149
transform 1 0 51980 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_559
timestamp 1644511149
transform 1 0 52532 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_561
timestamp 1644511149
transform 1 0 52716 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_573
timestamp 1644511149
transform 1 0 53820 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_585
timestamp 1644511149
transform 1 0 54924 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_597
timestamp 1644511149
transform 1 0 56028 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_609
timestamp 1644511149
transform 1 0 57132 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_615
timestamp 1644511149
transform 1 0 57684 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_65_617
timestamp 1644511149
transform 1 0 57868 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_66_3
timestamp 1644511149
transform 1 0 1380 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_15
timestamp 1644511149
transform 1 0 2484 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_66_27
timestamp 1644511149
transform 1 0 3588 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_29
timestamp 1644511149
transform 1 0 3772 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_41
timestamp 1644511149
transform 1 0 4876 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_53
timestamp 1644511149
transform 1 0 5980 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_65
timestamp 1644511149
transform 1 0 7084 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_77
timestamp 1644511149
transform 1 0 8188 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_83
timestamp 1644511149
transform 1 0 8740 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_85
timestamp 1644511149
transform 1 0 8924 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_97
timestamp 1644511149
transform 1 0 10028 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_109
timestamp 1644511149
transform 1 0 11132 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_121
timestamp 1644511149
transform 1 0 12236 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_133
timestamp 1644511149
transform 1 0 13340 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_139
timestamp 1644511149
transform 1 0 13892 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_141
timestamp 1644511149
transform 1 0 14076 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_153
timestamp 1644511149
transform 1 0 15180 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_165
timestamp 1644511149
transform 1 0 16284 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_177
timestamp 1644511149
transform 1 0 17388 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_189
timestamp 1644511149
transform 1 0 18492 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_195
timestamp 1644511149
transform 1 0 19044 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_197
timestamp 1644511149
transform 1 0 19228 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_209
timestamp 1644511149
transform 1 0 20332 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_221
timestamp 1644511149
transform 1 0 21436 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_233
timestamp 1644511149
transform 1 0 22540 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_245
timestamp 1644511149
transform 1 0 23644 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_251
timestamp 1644511149
transform 1 0 24196 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_253
timestamp 1644511149
transform 1 0 24380 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_265
timestamp 1644511149
transform 1 0 25484 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_277
timestamp 1644511149
transform 1 0 26588 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_289
timestamp 1644511149
transform 1 0 27692 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_301
timestamp 1644511149
transform 1 0 28796 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_307
timestamp 1644511149
transform 1 0 29348 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_309
timestamp 1644511149
transform 1 0 29532 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_321
timestamp 1644511149
transform 1 0 30636 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_333
timestamp 1644511149
transform 1 0 31740 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_345
timestamp 1644511149
transform 1 0 32844 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_357
timestamp 1644511149
transform 1 0 33948 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_363
timestamp 1644511149
transform 1 0 34500 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_365
timestamp 1644511149
transform 1 0 34684 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_377
timestamp 1644511149
transform 1 0 35788 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_389
timestamp 1644511149
transform 1 0 36892 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_401
timestamp 1644511149
transform 1 0 37996 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_413
timestamp 1644511149
transform 1 0 39100 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_419
timestamp 1644511149
transform 1 0 39652 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_421
timestamp 1644511149
transform 1 0 39836 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_433
timestamp 1644511149
transform 1 0 40940 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_445
timestamp 1644511149
transform 1 0 42044 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_457
timestamp 1644511149
transform 1 0 43148 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_469
timestamp 1644511149
transform 1 0 44252 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_475
timestamp 1644511149
transform 1 0 44804 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_477
timestamp 1644511149
transform 1 0 44988 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_489
timestamp 1644511149
transform 1 0 46092 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_501
timestamp 1644511149
transform 1 0 47196 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_513
timestamp 1644511149
transform 1 0 48300 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_525
timestamp 1644511149
transform 1 0 49404 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_531
timestamp 1644511149
transform 1 0 49956 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_533
timestamp 1644511149
transform 1 0 50140 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_545
timestamp 1644511149
transform 1 0 51244 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_557
timestamp 1644511149
transform 1 0 52348 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_569
timestamp 1644511149
transform 1 0 53452 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_581
timestamp 1644511149
transform 1 0 54556 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_587
timestamp 1644511149
transform 1 0 55108 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_589
timestamp 1644511149
transform 1 0 55292 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_601
timestamp 1644511149
transform 1 0 56396 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_613
timestamp 1644511149
transform 1 0 57500 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_3
timestamp 1644511149
transform 1 0 1380 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_15
timestamp 1644511149
transform 1 0 2484 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_27
timestamp 1644511149
transform 1 0 3588 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_39
timestamp 1644511149
transform 1 0 4692 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_67_51
timestamp 1644511149
transform 1 0 5796 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_67_55
timestamp 1644511149
transform 1 0 6164 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_57
timestamp 1644511149
transform 1 0 6348 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_69
timestamp 1644511149
transform 1 0 7452 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_81
timestamp 1644511149
transform 1 0 8556 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_93
timestamp 1644511149
transform 1 0 9660 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_105
timestamp 1644511149
transform 1 0 10764 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_111
timestamp 1644511149
transform 1 0 11316 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_113
timestamp 1644511149
transform 1 0 11500 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_125
timestamp 1644511149
transform 1 0 12604 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_137
timestamp 1644511149
transform 1 0 13708 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_149
timestamp 1644511149
transform 1 0 14812 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_161
timestamp 1644511149
transform 1 0 15916 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_167
timestamp 1644511149
transform 1 0 16468 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_169
timestamp 1644511149
transform 1 0 16652 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_181
timestamp 1644511149
transform 1 0 17756 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_193
timestamp 1644511149
transform 1 0 18860 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_205
timestamp 1644511149
transform 1 0 19964 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_217
timestamp 1644511149
transform 1 0 21068 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_223
timestamp 1644511149
transform 1 0 21620 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_225
timestamp 1644511149
transform 1 0 21804 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_237
timestamp 1644511149
transform 1 0 22908 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_249
timestamp 1644511149
transform 1 0 24012 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_261
timestamp 1644511149
transform 1 0 25116 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_273
timestamp 1644511149
transform 1 0 26220 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_279
timestamp 1644511149
transform 1 0 26772 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_281
timestamp 1644511149
transform 1 0 26956 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_293
timestamp 1644511149
transform 1 0 28060 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_305
timestamp 1644511149
transform 1 0 29164 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_317
timestamp 1644511149
transform 1 0 30268 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_329
timestamp 1644511149
transform 1 0 31372 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_335
timestamp 1644511149
transform 1 0 31924 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_337
timestamp 1644511149
transform 1 0 32108 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_349
timestamp 1644511149
transform 1 0 33212 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_361
timestamp 1644511149
transform 1 0 34316 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_373
timestamp 1644511149
transform 1 0 35420 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_385
timestamp 1644511149
transform 1 0 36524 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_391
timestamp 1644511149
transform 1 0 37076 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_393
timestamp 1644511149
transform 1 0 37260 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_405
timestamp 1644511149
transform 1 0 38364 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_417
timestamp 1644511149
transform 1 0 39468 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_429
timestamp 1644511149
transform 1 0 40572 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_441
timestamp 1644511149
transform 1 0 41676 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_447
timestamp 1644511149
transform 1 0 42228 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_449
timestamp 1644511149
transform 1 0 42412 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_461
timestamp 1644511149
transform 1 0 43516 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_473
timestamp 1644511149
transform 1 0 44620 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_485
timestamp 1644511149
transform 1 0 45724 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_497
timestamp 1644511149
transform 1 0 46828 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_503
timestamp 1644511149
transform 1 0 47380 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_505
timestamp 1644511149
transform 1 0 47564 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_517
timestamp 1644511149
transform 1 0 48668 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_529
timestamp 1644511149
transform 1 0 49772 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_541
timestamp 1644511149
transform 1 0 50876 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_553
timestamp 1644511149
transform 1 0 51980 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_559
timestamp 1644511149
transform 1 0 52532 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_561
timestamp 1644511149
transform 1 0 52716 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_573
timestamp 1644511149
transform 1 0 53820 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_585
timestamp 1644511149
transform 1 0 54924 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_597
timestamp 1644511149
transform 1 0 56028 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_609
timestamp 1644511149
transform 1 0 57132 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_615
timestamp 1644511149
transform 1 0 57684 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_67_617
timestamp 1644511149
transform 1 0 57868 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_68_3
timestamp 1644511149
transform 1 0 1380 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_15
timestamp 1644511149
transform 1 0 2484 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_68_27
timestamp 1644511149
transform 1 0 3588 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_29
timestamp 1644511149
transform 1 0 3772 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_41
timestamp 1644511149
transform 1 0 4876 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_53
timestamp 1644511149
transform 1 0 5980 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_65
timestamp 1644511149
transform 1 0 7084 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_77
timestamp 1644511149
transform 1 0 8188 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_83
timestamp 1644511149
transform 1 0 8740 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_85
timestamp 1644511149
transform 1 0 8924 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_97
timestamp 1644511149
transform 1 0 10028 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_109
timestamp 1644511149
transform 1 0 11132 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_121
timestamp 1644511149
transform 1 0 12236 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_133
timestamp 1644511149
transform 1 0 13340 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_139
timestamp 1644511149
transform 1 0 13892 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_141
timestamp 1644511149
transform 1 0 14076 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_153
timestamp 1644511149
transform 1 0 15180 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_165
timestamp 1644511149
transform 1 0 16284 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_177
timestamp 1644511149
transform 1 0 17388 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_189
timestamp 1644511149
transform 1 0 18492 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_195
timestamp 1644511149
transform 1 0 19044 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_197
timestamp 1644511149
transform 1 0 19228 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_209
timestamp 1644511149
transform 1 0 20332 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_221
timestamp 1644511149
transform 1 0 21436 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_233
timestamp 1644511149
transform 1 0 22540 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_245
timestamp 1644511149
transform 1 0 23644 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_251
timestamp 1644511149
transform 1 0 24196 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_253
timestamp 1644511149
transform 1 0 24380 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_265
timestamp 1644511149
transform 1 0 25484 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_277
timestamp 1644511149
transform 1 0 26588 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_289
timestamp 1644511149
transform 1 0 27692 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_301
timestamp 1644511149
transform 1 0 28796 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_307
timestamp 1644511149
transform 1 0 29348 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_309
timestamp 1644511149
transform 1 0 29532 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_321
timestamp 1644511149
transform 1 0 30636 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_333
timestamp 1644511149
transform 1 0 31740 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_345
timestamp 1644511149
transform 1 0 32844 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_357
timestamp 1644511149
transform 1 0 33948 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_363
timestamp 1644511149
transform 1 0 34500 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_365
timestamp 1644511149
transform 1 0 34684 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_377
timestamp 1644511149
transform 1 0 35788 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_389
timestamp 1644511149
transform 1 0 36892 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_401
timestamp 1644511149
transform 1 0 37996 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_413
timestamp 1644511149
transform 1 0 39100 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_419
timestamp 1644511149
transform 1 0 39652 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_421
timestamp 1644511149
transform 1 0 39836 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_433
timestamp 1644511149
transform 1 0 40940 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_445
timestamp 1644511149
transform 1 0 42044 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_457
timestamp 1644511149
transform 1 0 43148 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_469
timestamp 1644511149
transform 1 0 44252 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_475
timestamp 1644511149
transform 1 0 44804 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_477
timestamp 1644511149
transform 1 0 44988 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_489
timestamp 1644511149
transform 1 0 46092 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_501
timestamp 1644511149
transform 1 0 47196 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_513
timestamp 1644511149
transform 1 0 48300 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_525
timestamp 1644511149
transform 1 0 49404 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_531
timestamp 1644511149
transform 1 0 49956 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_533
timestamp 1644511149
transform 1 0 50140 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_545
timestamp 1644511149
transform 1 0 51244 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_557
timestamp 1644511149
transform 1 0 52348 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_569
timestamp 1644511149
transform 1 0 53452 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_581
timestamp 1644511149
transform 1 0 54556 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_587
timestamp 1644511149
transform 1 0 55108 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_589
timestamp 1644511149
transform 1 0 55292 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_601
timestamp 1644511149
transform 1 0 56396 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_613
timestamp 1644511149
transform 1 0 57500 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_3
timestamp 1644511149
transform 1 0 1380 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_15
timestamp 1644511149
transform 1 0 2484 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_27
timestamp 1644511149
transform 1 0 3588 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_39
timestamp 1644511149
transform 1 0 4692 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_69_51
timestamp 1644511149
transform 1 0 5796 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_69_55
timestamp 1644511149
transform 1 0 6164 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_57
timestamp 1644511149
transform 1 0 6348 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_69
timestamp 1644511149
transform 1 0 7452 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_81
timestamp 1644511149
transform 1 0 8556 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_93
timestamp 1644511149
transform 1 0 9660 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_105
timestamp 1644511149
transform 1 0 10764 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_111
timestamp 1644511149
transform 1 0 11316 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_113
timestamp 1644511149
transform 1 0 11500 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_125
timestamp 1644511149
transform 1 0 12604 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_137
timestamp 1644511149
transform 1 0 13708 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_149
timestamp 1644511149
transform 1 0 14812 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_161
timestamp 1644511149
transform 1 0 15916 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_167
timestamp 1644511149
transform 1 0 16468 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_169
timestamp 1644511149
transform 1 0 16652 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_181
timestamp 1644511149
transform 1 0 17756 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_193
timestamp 1644511149
transform 1 0 18860 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_205
timestamp 1644511149
transform 1 0 19964 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_217
timestamp 1644511149
transform 1 0 21068 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_223
timestamp 1644511149
transform 1 0 21620 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_225
timestamp 1644511149
transform 1 0 21804 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_237
timestamp 1644511149
transform 1 0 22908 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_249
timestamp 1644511149
transform 1 0 24012 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_261
timestamp 1644511149
transform 1 0 25116 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_273
timestamp 1644511149
transform 1 0 26220 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_279
timestamp 1644511149
transform 1 0 26772 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_281
timestamp 1644511149
transform 1 0 26956 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_293
timestamp 1644511149
transform 1 0 28060 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_305
timestamp 1644511149
transform 1 0 29164 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_317
timestamp 1644511149
transform 1 0 30268 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_329
timestamp 1644511149
transform 1 0 31372 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_335
timestamp 1644511149
transform 1 0 31924 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_337
timestamp 1644511149
transform 1 0 32108 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_349
timestamp 1644511149
transform 1 0 33212 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_361
timestamp 1644511149
transform 1 0 34316 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_373
timestamp 1644511149
transform 1 0 35420 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_385
timestamp 1644511149
transform 1 0 36524 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_391
timestamp 1644511149
transform 1 0 37076 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_393
timestamp 1644511149
transform 1 0 37260 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_405
timestamp 1644511149
transform 1 0 38364 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_417
timestamp 1644511149
transform 1 0 39468 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_429
timestamp 1644511149
transform 1 0 40572 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_441
timestamp 1644511149
transform 1 0 41676 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_447
timestamp 1644511149
transform 1 0 42228 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_449
timestamp 1644511149
transform 1 0 42412 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_461
timestamp 1644511149
transform 1 0 43516 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_473
timestamp 1644511149
transform 1 0 44620 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_485
timestamp 1644511149
transform 1 0 45724 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_497
timestamp 1644511149
transform 1 0 46828 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_503
timestamp 1644511149
transform 1 0 47380 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_505
timestamp 1644511149
transform 1 0 47564 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_517
timestamp 1644511149
transform 1 0 48668 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_529
timestamp 1644511149
transform 1 0 49772 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_541
timestamp 1644511149
transform 1 0 50876 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_553
timestamp 1644511149
transform 1 0 51980 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_559
timestamp 1644511149
transform 1 0 52532 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_561
timestamp 1644511149
transform 1 0 52716 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_573
timestamp 1644511149
transform 1 0 53820 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_585
timestamp 1644511149
transform 1 0 54924 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_597
timestamp 1644511149
transform 1 0 56028 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_609
timestamp 1644511149
transform 1 0 57132 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_615
timestamp 1644511149
transform 1 0 57684 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_69_617
timestamp 1644511149
transform 1 0 57868 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_70_3
timestamp 1644511149
transform 1 0 1380 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_15
timestamp 1644511149
transform 1 0 2484 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_70_27
timestamp 1644511149
transform 1 0 3588 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_29
timestamp 1644511149
transform 1 0 3772 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_41
timestamp 1644511149
transform 1 0 4876 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_53
timestamp 1644511149
transform 1 0 5980 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_65
timestamp 1644511149
transform 1 0 7084 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_77
timestamp 1644511149
transform 1 0 8188 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_83
timestamp 1644511149
transform 1 0 8740 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_85
timestamp 1644511149
transform 1 0 8924 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_97
timestamp 1644511149
transform 1 0 10028 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_109
timestamp 1644511149
transform 1 0 11132 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_121
timestamp 1644511149
transform 1 0 12236 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_133
timestamp 1644511149
transform 1 0 13340 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_139
timestamp 1644511149
transform 1 0 13892 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_141
timestamp 1644511149
transform 1 0 14076 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_153
timestamp 1644511149
transform 1 0 15180 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_165
timestamp 1644511149
transform 1 0 16284 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_177
timestamp 1644511149
transform 1 0 17388 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_189
timestamp 1644511149
transform 1 0 18492 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_195
timestamp 1644511149
transform 1 0 19044 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_197
timestamp 1644511149
transform 1 0 19228 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_209
timestamp 1644511149
transform 1 0 20332 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_221
timestamp 1644511149
transform 1 0 21436 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_233
timestamp 1644511149
transform 1 0 22540 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_245
timestamp 1644511149
transform 1 0 23644 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_251
timestamp 1644511149
transform 1 0 24196 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_253
timestamp 1644511149
transform 1 0 24380 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_265
timestamp 1644511149
transform 1 0 25484 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_277
timestamp 1644511149
transform 1 0 26588 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_289
timestamp 1644511149
transform 1 0 27692 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_301
timestamp 1644511149
transform 1 0 28796 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_307
timestamp 1644511149
transform 1 0 29348 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_309
timestamp 1644511149
transform 1 0 29532 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_321
timestamp 1644511149
transform 1 0 30636 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_333
timestamp 1644511149
transform 1 0 31740 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_345
timestamp 1644511149
transform 1 0 32844 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_357
timestamp 1644511149
transform 1 0 33948 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_363
timestamp 1644511149
transform 1 0 34500 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_365
timestamp 1644511149
transform 1 0 34684 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_377
timestamp 1644511149
transform 1 0 35788 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_389
timestamp 1644511149
transform 1 0 36892 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_401
timestamp 1644511149
transform 1 0 37996 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_413
timestamp 1644511149
transform 1 0 39100 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_419
timestamp 1644511149
transform 1 0 39652 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_421
timestamp 1644511149
transform 1 0 39836 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_433
timestamp 1644511149
transform 1 0 40940 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_445
timestamp 1644511149
transform 1 0 42044 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_457
timestamp 1644511149
transform 1 0 43148 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_469
timestamp 1644511149
transform 1 0 44252 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_475
timestamp 1644511149
transform 1 0 44804 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_477
timestamp 1644511149
transform 1 0 44988 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_489
timestamp 1644511149
transform 1 0 46092 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_501
timestamp 1644511149
transform 1 0 47196 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_513
timestamp 1644511149
transform 1 0 48300 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_525
timestamp 1644511149
transform 1 0 49404 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_531
timestamp 1644511149
transform 1 0 49956 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_533
timestamp 1644511149
transform 1 0 50140 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_545
timestamp 1644511149
transform 1 0 51244 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_557
timestamp 1644511149
transform 1 0 52348 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_569
timestamp 1644511149
transform 1 0 53452 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_581
timestamp 1644511149
transform 1 0 54556 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_587
timestamp 1644511149
transform 1 0 55108 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_589
timestamp 1644511149
transform 1 0 55292 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_601
timestamp 1644511149
transform 1 0 56396 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_613
timestamp 1644511149
transform 1 0 57500 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_3
timestamp 1644511149
transform 1 0 1380 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_15
timestamp 1644511149
transform 1 0 2484 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_27
timestamp 1644511149
transform 1 0 3588 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_39
timestamp 1644511149
transform 1 0 4692 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_71_51
timestamp 1644511149
transform 1 0 5796 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_71_55
timestamp 1644511149
transform 1 0 6164 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_57
timestamp 1644511149
transform 1 0 6348 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_69
timestamp 1644511149
transform 1 0 7452 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_81
timestamp 1644511149
transform 1 0 8556 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_93
timestamp 1644511149
transform 1 0 9660 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_105
timestamp 1644511149
transform 1 0 10764 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_111
timestamp 1644511149
transform 1 0 11316 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_113
timestamp 1644511149
transform 1 0 11500 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_125
timestamp 1644511149
transform 1 0 12604 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_137
timestamp 1644511149
transform 1 0 13708 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_149
timestamp 1644511149
transform 1 0 14812 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_161
timestamp 1644511149
transform 1 0 15916 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_167
timestamp 1644511149
transform 1 0 16468 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_169
timestamp 1644511149
transform 1 0 16652 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_181
timestamp 1644511149
transform 1 0 17756 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_193
timestamp 1644511149
transform 1 0 18860 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_205
timestamp 1644511149
transform 1 0 19964 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_217
timestamp 1644511149
transform 1 0 21068 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_223
timestamp 1644511149
transform 1 0 21620 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_225
timestamp 1644511149
transform 1 0 21804 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_237
timestamp 1644511149
transform 1 0 22908 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_249
timestamp 1644511149
transform 1 0 24012 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_261
timestamp 1644511149
transform 1 0 25116 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_273
timestamp 1644511149
transform 1 0 26220 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_279
timestamp 1644511149
transform 1 0 26772 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_281
timestamp 1644511149
transform 1 0 26956 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_293
timestamp 1644511149
transform 1 0 28060 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_305
timestamp 1644511149
transform 1 0 29164 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_317
timestamp 1644511149
transform 1 0 30268 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_329
timestamp 1644511149
transform 1 0 31372 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_335
timestamp 1644511149
transform 1 0 31924 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_337
timestamp 1644511149
transform 1 0 32108 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_349
timestamp 1644511149
transform 1 0 33212 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_361
timestamp 1644511149
transform 1 0 34316 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_373
timestamp 1644511149
transform 1 0 35420 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_385
timestamp 1644511149
transform 1 0 36524 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_391
timestamp 1644511149
transform 1 0 37076 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_393
timestamp 1644511149
transform 1 0 37260 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_405
timestamp 1644511149
transform 1 0 38364 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_417
timestamp 1644511149
transform 1 0 39468 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_429
timestamp 1644511149
transform 1 0 40572 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_441
timestamp 1644511149
transform 1 0 41676 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_447
timestamp 1644511149
transform 1 0 42228 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_449
timestamp 1644511149
transform 1 0 42412 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_461
timestamp 1644511149
transform 1 0 43516 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_71_473
timestamp 1644511149
transform 1 0 44620 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_71_481
timestamp 1644511149
transform 1 0 45356 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_71_486
timestamp 1644511149
transform 1 0 45816 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_498
timestamp 1644511149
transform 1 0 46920 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_71_505
timestamp 1644511149
transform 1 0 47564 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_517
timestamp 1644511149
transform 1 0 48668 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_529
timestamp 1644511149
transform 1 0 49772 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_541
timestamp 1644511149
transform 1 0 50876 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_553
timestamp 1644511149
transform 1 0 51980 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_559
timestamp 1644511149
transform 1 0 52532 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_561
timestamp 1644511149
transform 1 0 52716 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_573
timestamp 1644511149
transform 1 0 53820 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_585
timestamp 1644511149
transform 1 0 54924 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_597
timestamp 1644511149
transform 1 0 56028 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_609
timestamp 1644511149
transform 1 0 57132 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_615
timestamp 1644511149
transform 1 0 57684 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_71_617
timestamp 1644511149
transform 1 0 57868 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_72_3
timestamp 1644511149
transform 1 0 1380 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_15
timestamp 1644511149
transform 1 0 2484 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_72_27
timestamp 1644511149
transform 1 0 3588 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_29
timestamp 1644511149
transform 1 0 3772 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_41
timestamp 1644511149
transform 1 0 4876 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_53
timestamp 1644511149
transform 1 0 5980 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_65
timestamp 1644511149
transform 1 0 7084 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_77
timestamp 1644511149
transform 1 0 8188 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_83
timestamp 1644511149
transform 1 0 8740 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_85
timestamp 1644511149
transform 1 0 8924 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_97
timestamp 1644511149
transform 1 0 10028 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_109
timestamp 1644511149
transform 1 0 11132 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_121
timestamp 1644511149
transform 1 0 12236 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_133
timestamp 1644511149
transform 1 0 13340 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_139
timestamp 1644511149
transform 1 0 13892 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_141
timestamp 1644511149
transform 1 0 14076 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_153
timestamp 1644511149
transform 1 0 15180 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_165
timestamp 1644511149
transform 1 0 16284 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_177
timestamp 1644511149
transform 1 0 17388 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_189
timestamp 1644511149
transform 1 0 18492 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_195
timestamp 1644511149
transform 1 0 19044 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_197
timestamp 1644511149
transform 1 0 19228 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_209
timestamp 1644511149
transform 1 0 20332 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_221
timestamp 1644511149
transform 1 0 21436 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_233
timestamp 1644511149
transform 1 0 22540 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_245
timestamp 1644511149
transform 1 0 23644 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_251
timestamp 1644511149
transform 1 0 24196 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_253
timestamp 1644511149
transform 1 0 24380 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_265
timestamp 1644511149
transform 1 0 25484 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_277
timestamp 1644511149
transform 1 0 26588 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_289
timestamp 1644511149
transform 1 0 27692 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_301
timestamp 1644511149
transform 1 0 28796 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_307
timestamp 1644511149
transform 1 0 29348 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_309
timestamp 1644511149
transform 1 0 29532 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_321
timestamp 1644511149
transform 1 0 30636 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_333
timestamp 1644511149
transform 1 0 31740 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_345
timestamp 1644511149
transform 1 0 32844 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_357
timestamp 1644511149
transform 1 0 33948 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_363
timestamp 1644511149
transform 1 0 34500 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_365
timestamp 1644511149
transform 1 0 34684 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_377
timestamp 1644511149
transform 1 0 35788 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_389
timestamp 1644511149
transform 1 0 36892 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_401
timestamp 1644511149
transform 1 0 37996 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_413
timestamp 1644511149
transform 1 0 39100 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_419
timestamp 1644511149
transform 1 0 39652 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_421
timestamp 1644511149
transform 1 0 39836 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_433
timestamp 1644511149
transform 1 0 40940 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_445
timestamp 1644511149
transform 1 0 42044 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_457
timestamp 1644511149
transform 1 0 43148 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_469
timestamp 1644511149
transform 1 0 44252 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_475
timestamp 1644511149
transform 1 0 44804 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_72_480
timestamp 1644511149
transform 1 0 45264 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_72_484
timestamp 1644511149
transform 1 0 45632 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_501
timestamp 1644511149
transform 1 0 47196 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_513
timestamp 1644511149
transform 1 0 48300 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_525
timestamp 1644511149
transform 1 0 49404 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_531
timestamp 1644511149
transform 1 0 49956 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_533
timestamp 1644511149
transform 1 0 50140 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_72_545
timestamp 1644511149
transform 1 0 51244 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_72_549
timestamp 1644511149
transform 1 0 51612 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_562
timestamp 1644511149
transform 1 0 52808 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_574
timestamp 1644511149
transform 1 0 53912 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_72_586
timestamp 1644511149
transform 1 0 55016 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_72_589
timestamp 1644511149
transform 1 0 55292 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_72_597
timestamp 1644511149
transform 1 0 56028 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_72_621
timestamp 1644511149
transform 1 0 58236 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_73_3
timestamp 1644511149
transform 1 0 1380 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_73_11
timestamp 1644511149
transform 1 0 2116 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_73_34
timestamp 1644511149
transform 1 0 4232 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_73_46
timestamp 1644511149
transform 1 0 5336 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_73_54
timestamp 1644511149
transform 1 0 6072 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_73_57
timestamp 1644511149
transform 1 0 6348 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_69
timestamp 1644511149
transform 1 0 7452 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_81
timestamp 1644511149
transform 1 0 8556 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_93
timestamp 1644511149
transform 1 0 9660 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_105
timestamp 1644511149
transform 1 0 10764 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_111
timestamp 1644511149
transform 1 0 11316 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_113
timestamp 1644511149
transform 1 0 11500 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_125
timestamp 1644511149
transform 1 0 12604 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_137
timestamp 1644511149
transform 1 0 13708 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_149
timestamp 1644511149
transform 1 0 14812 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_161
timestamp 1644511149
transform 1 0 15916 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_167
timestamp 1644511149
transform 1 0 16468 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_169
timestamp 1644511149
transform 1 0 16652 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_181
timestamp 1644511149
transform 1 0 17756 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_193
timestamp 1644511149
transform 1 0 18860 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_205
timestamp 1644511149
transform 1 0 19964 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_217
timestamp 1644511149
transform 1 0 21068 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_223
timestamp 1644511149
transform 1 0 21620 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_225
timestamp 1644511149
transform 1 0 21804 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_237
timestamp 1644511149
transform 1 0 22908 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_249
timestamp 1644511149
transform 1 0 24012 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_261
timestamp 1644511149
transform 1 0 25116 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_273
timestamp 1644511149
transform 1 0 26220 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_279
timestamp 1644511149
transform 1 0 26772 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_281
timestamp 1644511149
transform 1 0 26956 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_293
timestamp 1644511149
transform 1 0 28060 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_305
timestamp 1644511149
transform 1 0 29164 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_317
timestamp 1644511149
transform 1 0 30268 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_329
timestamp 1644511149
transform 1 0 31372 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_335
timestamp 1644511149
transform 1 0 31924 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_337
timestamp 1644511149
transform 1 0 32108 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_349
timestamp 1644511149
transform 1 0 33212 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_361
timestamp 1644511149
transform 1 0 34316 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_373
timestamp 1644511149
transform 1 0 35420 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_385
timestamp 1644511149
transform 1 0 36524 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_391
timestamp 1644511149
transform 1 0 37076 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_393
timestamp 1644511149
transform 1 0 37260 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_405
timestamp 1644511149
transform 1 0 38364 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_417
timestamp 1644511149
transform 1 0 39468 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_429
timestamp 1644511149
transform 1 0 40572 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_441
timestamp 1644511149
transform 1 0 41676 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_447
timestamp 1644511149
transform 1 0 42228 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_449
timestamp 1644511149
transform 1 0 42412 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_73_461
timestamp 1644511149
transform 1 0 43516 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_73_465
timestamp 1644511149
transform 1 0 43884 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_73_470
timestamp 1644511149
transform 1 0 44344 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_73_474
timestamp 1644511149
transform 1 0 44712 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_73_479
timestamp 1644511149
transform 1 0 45172 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_73_499
timestamp 1644511149
transform 1 0 47012 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_73_503
timestamp 1644511149
transform 1 0 47380 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_73_505
timestamp 1644511149
transform 1 0 47564 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_73_513
timestamp 1644511149
transform 1 0 48300 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_73_535
timestamp 1644511149
transform 1 0 50324 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_73_555
timestamp 1644511149
transform 1 0 52164 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_73_559
timestamp 1644511149
transform 1 0 52532 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_573
timestamp 1644511149
transform 1 0 53820 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_585
timestamp 1644511149
transform 1 0 54924 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_597
timestamp 1644511149
transform 1 0 56028 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_603
timestamp 1644511149
transform 1 0 56580 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_73_607
timestamp 1644511149
transform 1 0 56948 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_73_615
timestamp 1644511149
transform 1 0 57684 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_73_617
timestamp 1644511149
transform 1 0 57868 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_74_3
timestamp 1644511149
transform 1 0 1380 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_15
timestamp 1644511149
transform 1 0 2484 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_74_27
timestamp 1644511149
transform 1 0 3588 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_32
timestamp 1644511149
transform 1 0 4048 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_44
timestamp 1644511149
transform 1 0 5152 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_56
timestamp 1644511149
transform 1 0 6256 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_68
timestamp 1644511149
transform 1 0 7360 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_74_80
timestamp 1644511149
transform 1 0 8464 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_74_85
timestamp 1644511149
transform 1 0 8924 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_97
timestamp 1644511149
transform 1 0 10028 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_109
timestamp 1644511149
transform 1 0 11132 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_121
timestamp 1644511149
transform 1 0 12236 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_133
timestamp 1644511149
transform 1 0 13340 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_139
timestamp 1644511149
transform 1 0 13892 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_141
timestamp 1644511149
transform 1 0 14076 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_153
timestamp 1644511149
transform 1 0 15180 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_165
timestamp 1644511149
transform 1 0 16284 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_177
timestamp 1644511149
transform 1 0 17388 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_189
timestamp 1644511149
transform 1 0 18492 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_195
timestamp 1644511149
transform 1 0 19044 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_197
timestamp 1644511149
transform 1 0 19228 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_209
timestamp 1644511149
transform 1 0 20332 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_221
timestamp 1644511149
transform 1 0 21436 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_233
timestamp 1644511149
transform 1 0 22540 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_245
timestamp 1644511149
transform 1 0 23644 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_251
timestamp 1644511149
transform 1 0 24196 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_253
timestamp 1644511149
transform 1 0 24380 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_265
timestamp 1644511149
transform 1 0 25484 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_277
timestamp 1644511149
transform 1 0 26588 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_289
timestamp 1644511149
transform 1 0 27692 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_301
timestamp 1644511149
transform 1 0 28796 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_307
timestamp 1644511149
transform 1 0 29348 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_309
timestamp 1644511149
transform 1 0 29532 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_321
timestamp 1644511149
transform 1 0 30636 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_333
timestamp 1644511149
transform 1 0 31740 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_345
timestamp 1644511149
transform 1 0 32844 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_357
timestamp 1644511149
transform 1 0 33948 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_363
timestamp 1644511149
transform 1 0 34500 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_365
timestamp 1644511149
transform 1 0 34684 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_74_377
timestamp 1644511149
transform 1 0 35788 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_74_385
timestamp 1644511149
transform 1 0 36524 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_402
timestamp 1644511149
transform 1 0 38088 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_414
timestamp 1644511149
transform 1 0 39192 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_74_421
timestamp 1644511149
transform 1 0 39836 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_74_444
timestamp 1644511149
transform 1 0 41952 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_74_472
timestamp 1644511149
transform 1 0 44528 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_74_482
timestamp 1644511149
transform 1 0 45448 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_74_490
timestamp 1644511149
transform 1 0 46184 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_74_502
timestamp 1644511149
transform 1 0 47288 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_74_506
timestamp 1644511149
transform 1 0 47656 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_74_528
timestamp 1644511149
transform 1 0 49680 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_74_533
timestamp 1644511149
transform 1 0 50140 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_74_547
timestamp 1644511149
transform 1 0 51428 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_74_572
timestamp 1644511149
transform 1 0 53728 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_74_584
timestamp 1644511149
transform 1 0 54832 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_74_589
timestamp 1644511149
transform 1 0 55292 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_74_601
timestamp 1644511149
transform 1 0 56396 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_74_609
timestamp 1644511149
transform 1 0 57132 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_613
timestamp 1644511149
transform 1 0 57500 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_75_3
timestamp 1644511149
transform 1 0 1380 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_75_11
timestamp 1644511149
transform 1 0 2116 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_75_17
timestamp 1644511149
transform 1 0 2668 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_29
timestamp 1644511149
transform 1 0 3772 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_41
timestamp 1644511149
transform 1 0 4876 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_75_53
timestamp 1644511149
transform 1 0 5980 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_75_57
timestamp 1644511149
transform 1 0 6348 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_69
timestamp 1644511149
transform 1 0 7452 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_81
timestamp 1644511149
transform 1 0 8556 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_93
timestamp 1644511149
transform 1 0 9660 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_105
timestamp 1644511149
transform 1 0 10764 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_111
timestamp 1644511149
transform 1 0 11316 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_113
timestamp 1644511149
transform 1 0 11500 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_125
timestamp 1644511149
transform 1 0 12604 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_137
timestamp 1644511149
transform 1 0 13708 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_149
timestamp 1644511149
transform 1 0 14812 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_161
timestamp 1644511149
transform 1 0 15916 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_167
timestamp 1644511149
transform 1 0 16468 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_169
timestamp 1644511149
transform 1 0 16652 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_181
timestamp 1644511149
transform 1 0 17756 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_193
timestamp 1644511149
transform 1 0 18860 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_205
timestamp 1644511149
transform 1 0 19964 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_217
timestamp 1644511149
transform 1 0 21068 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_223
timestamp 1644511149
transform 1 0 21620 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_225
timestamp 1644511149
transform 1 0 21804 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_237
timestamp 1644511149
transform 1 0 22908 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_249
timestamp 1644511149
transform 1 0 24012 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_261
timestamp 1644511149
transform 1 0 25116 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_273
timestamp 1644511149
transform 1 0 26220 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_279
timestamp 1644511149
transform 1 0 26772 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_281
timestamp 1644511149
transform 1 0 26956 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_293
timestamp 1644511149
transform 1 0 28060 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_305
timestamp 1644511149
transform 1 0 29164 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_317
timestamp 1644511149
transform 1 0 30268 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_329
timestamp 1644511149
transform 1 0 31372 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_335
timestamp 1644511149
transform 1 0 31924 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_337
timestamp 1644511149
transform 1 0 32108 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_349
timestamp 1644511149
transform 1 0 33212 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_361
timestamp 1644511149
transform 1 0 34316 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_373
timestamp 1644511149
transform 1 0 35420 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_75_388
timestamp 1644511149
transform 1 0 36800 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_75_409
timestamp 1644511149
transform 1 0 38732 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_442
timestamp 1644511149
transform 1 0 41768 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_75_449
timestamp 1644511149
transform 1 0 42412 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_75_461
timestamp 1644511149
transform 1 0 43516 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_75_470
timestamp 1644511149
transform 1 0 44344 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_75_484
timestamp 1644511149
transform 1 0 45632 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_75_495
timestamp 1644511149
transform 1 0 46644 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_75_503
timestamp 1644511149
transform 1 0 47380 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_75_505
timestamp 1644511149
transform 1 0 47564 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_511
timestamp 1644511149
transform 1 0 48116 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_533
timestamp 1644511149
transform 1 0 50140 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_545
timestamp 1644511149
transform 1 0 51244 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_75_557
timestamp 1644511149
transform 1 0 52348 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_75_567
timestamp 1644511149
transform 1 0 53268 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_579
timestamp 1644511149
transform 1 0 54372 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_591
timestamp 1644511149
transform 1 0 55476 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_603
timestamp 1644511149
transform 1 0 56580 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_75_615
timestamp 1644511149
transform 1 0 57684 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_75_617
timestamp 1644511149
transform 1 0 57868 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_76_3
timestamp 1644511149
transform 1 0 1380 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_15
timestamp 1644511149
transform 1 0 2484 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_76_27
timestamp 1644511149
transform 1 0 3588 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_29
timestamp 1644511149
transform 1 0 3772 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_41
timestamp 1644511149
transform 1 0 4876 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_53
timestamp 1644511149
transform 1 0 5980 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_65
timestamp 1644511149
transform 1 0 7084 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_77
timestamp 1644511149
transform 1 0 8188 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_83
timestamp 1644511149
transform 1 0 8740 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_85
timestamp 1644511149
transform 1 0 8924 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_97
timestamp 1644511149
transform 1 0 10028 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_109
timestamp 1644511149
transform 1 0 11132 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_121
timestamp 1644511149
transform 1 0 12236 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_133
timestamp 1644511149
transform 1 0 13340 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_139
timestamp 1644511149
transform 1 0 13892 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_141
timestamp 1644511149
transform 1 0 14076 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_153
timestamp 1644511149
transform 1 0 15180 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_165
timestamp 1644511149
transform 1 0 16284 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_177
timestamp 1644511149
transform 1 0 17388 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_189
timestamp 1644511149
transform 1 0 18492 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_195
timestamp 1644511149
transform 1 0 19044 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_197
timestamp 1644511149
transform 1 0 19228 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_209
timestamp 1644511149
transform 1 0 20332 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_221
timestamp 1644511149
transform 1 0 21436 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_233
timestamp 1644511149
transform 1 0 22540 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_245
timestamp 1644511149
transform 1 0 23644 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_251
timestamp 1644511149
transform 1 0 24196 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_253
timestamp 1644511149
transform 1 0 24380 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_265
timestamp 1644511149
transform 1 0 25484 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_277
timestamp 1644511149
transform 1 0 26588 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_289
timestamp 1644511149
transform 1 0 27692 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_301
timestamp 1644511149
transform 1 0 28796 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_307
timestamp 1644511149
transform 1 0 29348 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_309
timestamp 1644511149
transform 1 0 29532 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_321
timestamp 1644511149
transform 1 0 30636 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_333
timestamp 1644511149
transform 1 0 31740 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_345
timestamp 1644511149
transform 1 0 32844 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_357
timestamp 1644511149
transform 1 0 33948 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_363
timestamp 1644511149
transform 1 0 34500 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_365
timestamp 1644511149
transform 1 0 34684 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_377
timestamp 1644511149
transform 1 0 35788 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_76_389
timestamp 1644511149
transform 1 0 36892 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_76_397
timestamp 1644511149
transform 1 0 37628 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_76_405
timestamp 1644511149
transform 1 0 38364 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_76_417
timestamp 1644511149
transform 1 0 39468 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_76_421
timestamp 1644511149
transform 1 0 39836 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_427
timestamp 1644511149
transform 1 0 40388 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_440
timestamp 1644511149
transform 1 0 41584 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_452
timestamp 1644511149
transform 1 0 42688 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_76_464
timestamp 1644511149
transform 1 0 43792 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_76_470
timestamp 1644511149
transform 1 0 44344 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_76_477
timestamp 1644511149
transform 1 0 44988 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_76_489
timestamp 1644511149
transform 1 0 46092 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_76_493
timestamp 1644511149
transform 1 0 46460 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_497
timestamp 1644511149
transform 1 0 46828 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_509
timestamp 1644511149
transform 1 0 47932 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_76_521
timestamp 1644511149
transform 1 0 49036 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_76_529
timestamp 1644511149
transform 1 0 49772 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_76_533
timestamp 1644511149
transform 1 0 50140 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_545
timestamp 1644511149
transform 1 0 51244 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_557
timestamp 1644511149
transform 1 0 52348 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_569
timestamp 1644511149
transform 1 0 53452 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_581
timestamp 1644511149
transform 1 0 54556 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_587
timestamp 1644511149
transform 1 0 55108 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_589
timestamp 1644511149
transform 1 0 55292 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_601
timestamp 1644511149
transform 1 0 56396 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_613
timestamp 1644511149
transform 1 0 57500 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_3
timestamp 1644511149
transform 1 0 1380 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_77_30
timestamp 1644511149
transform 1 0 3864 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_42
timestamp 1644511149
transform 1 0 4968 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_77_54
timestamp 1644511149
transform 1 0 6072 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_77_57
timestamp 1644511149
transform 1 0 6348 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_69
timestamp 1644511149
transform 1 0 7452 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_81
timestamp 1644511149
transform 1 0 8556 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_93
timestamp 1644511149
transform 1 0 9660 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_105
timestamp 1644511149
transform 1 0 10764 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_111
timestamp 1644511149
transform 1 0 11316 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_113
timestamp 1644511149
transform 1 0 11500 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_125
timestamp 1644511149
transform 1 0 12604 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_137
timestamp 1644511149
transform 1 0 13708 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_149
timestamp 1644511149
transform 1 0 14812 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_161
timestamp 1644511149
transform 1 0 15916 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_167
timestamp 1644511149
transform 1 0 16468 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_169
timestamp 1644511149
transform 1 0 16652 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_181
timestamp 1644511149
transform 1 0 17756 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_193
timestamp 1644511149
transform 1 0 18860 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_205
timestamp 1644511149
transform 1 0 19964 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_217
timestamp 1644511149
transform 1 0 21068 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_223
timestamp 1644511149
transform 1 0 21620 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_225
timestamp 1644511149
transform 1 0 21804 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_237
timestamp 1644511149
transform 1 0 22908 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_249
timestamp 1644511149
transform 1 0 24012 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_261
timestamp 1644511149
transform 1 0 25116 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_273
timestamp 1644511149
transform 1 0 26220 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_279
timestamp 1644511149
transform 1 0 26772 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_281
timestamp 1644511149
transform 1 0 26956 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_293
timestamp 1644511149
transform 1 0 28060 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_305
timestamp 1644511149
transform 1 0 29164 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_317
timestamp 1644511149
transform 1 0 30268 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_329
timestamp 1644511149
transform 1 0 31372 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_335
timestamp 1644511149
transform 1 0 31924 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_337
timestamp 1644511149
transform 1 0 32108 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_349
timestamp 1644511149
transform 1 0 33212 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_361
timestamp 1644511149
transform 1 0 34316 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_373
timestamp 1644511149
transform 1 0 35420 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_385
timestamp 1644511149
transform 1 0 36524 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_391
timestamp 1644511149
transform 1 0 37076 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_77_409
timestamp 1644511149
transform 1 0 38732 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_77_420
timestamp 1644511149
transform 1 0 39744 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_77_436
timestamp 1644511149
transform 1 0 41216 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_449
timestamp 1644511149
transform 1 0 42412 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_77_461
timestamp 1644511149
transform 1 0 43516 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_77_466
timestamp 1644511149
transform 1 0 43976 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_472
timestamp 1644511149
transform 1 0 44528 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_77_483
timestamp 1644511149
transform 1 0 45540 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_489
timestamp 1644511149
transform 1 0 46092 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_77_494
timestamp 1644511149
transform 1 0 46552 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_77_502
timestamp 1644511149
transform 1 0 47288 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_77_505
timestamp 1644511149
transform 1 0 47564 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_77_517
timestamp 1644511149
transform 1 0 48668 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_77_521
timestamp 1644511149
transform 1 0 49036 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_543
timestamp 1644511149
transform 1 0 51060 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_77_555
timestamp 1644511149
transform 1 0 52164 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_77_559
timestamp 1644511149
transform 1 0 52532 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_565
timestamp 1644511149
transform 1 0 53084 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_577
timestamp 1644511149
transform 1 0 54188 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_589
timestamp 1644511149
transform 1 0 55292 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_601
timestamp 1644511149
transform 1 0 56396 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_77_613
timestamp 1644511149
transform 1 0 57500 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_77_617
timestamp 1644511149
transform 1 0 57868 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_78_3
timestamp 1644511149
transform 1 0 1380 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_78_11
timestamp 1644511149
transform 1 0 2116 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_78_16
timestamp 1644511149
transform 1 0 2576 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_29
timestamp 1644511149
transform 1 0 3772 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_41
timestamp 1644511149
transform 1 0 4876 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_53
timestamp 1644511149
transform 1 0 5980 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_65
timestamp 1644511149
transform 1 0 7084 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_77
timestamp 1644511149
transform 1 0 8188 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_83
timestamp 1644511149
transform 1 0 8740 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_85
timestamp 1644511149
transform 1 0 8924 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_97
timestamp 1644511149
transform 1 0 10028 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_109
timestamp 1644511149
transform 1 0 11132 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_121
timestamp 1644511149
transform 1 0 12236 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_133
timestamp 1644511149
transform 1 0 13340 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_139
timestamp 1644511149
transform 1 0 13892 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_141
timestamp 1644511149
transform 1 0 14076 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_153
timestamp 1644511149
transform 1 0 15180 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_165
timestamp 1644511149
transform 1 0 16284 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_177
timestamp 1644511149
transform 1 0 17388 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_189
timestamp 1644511149
transform 1 0 18492 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_195
timestamp 1644511149
transform 1 0 19044 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_197
timestamp 1644511149
transform 1 0 19228 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_209
timestamp 1644511149
transform 1 0 20332 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_221
timestamp 1644511149
transform 1 0 21436 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_233
timestamp 1644511149
transform 1 0 22540 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_245
timestamp 1644511149
transform 1 0 23644 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_251
timestamp 1644511149
transform 1 0 24196 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_253
timestamp 1644511149
transform 1 0 24380 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_265
timestamp 1644511149
transform 1 0 25484 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_277
timestamp 1644511149
transform 1 0 26588 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_289
timestamp 1644511149
transform 1 0 27692 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_301
timestamp 1644511149
transform 1 0 28796 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_307
timestamp 1644511149
transform 1 0 29348 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_309
timestamp 1644511149
transform 1 0 29532 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_321
timestamp 1644511149
transform 1 0 30636 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_333
timestamp 1644511149
transform 1 0 31740 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_345
timestamp 1644511149
transform 1 0 32844 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_357
timestamp 1644511149
transform 1 0 33948 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_363
timestamp 1644511149
transform 1 0 34500 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_365
timestamp 1644511149
transform 1 0 34684 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_78_377
timestamp 1644511149
transform 1 0 35788 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_78_385
timestamp 1644511149
transform 1 0 36524 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_78_391
timestamp 1644511149
transform 1 0 37076 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_78_399
timestamp 1644511149
transform 1 0 37812 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_78_411
timestamp 1644511149
transform 1 0 38916 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_78_419
timestamp 1644511149
transform 1 0 39652 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_442
timestamp 1644511149
transform 1 0 41768 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_78_454
timestamp 1644511149
transform 1 0 42872 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_78_472
timestamp 1644511149
transform 1 0 44528 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_78_477
timestamp 1644511149
transform 1 0 44988 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_78_487
timestamp 1644511149
transform 1 0 45908 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_78_499
timestamp 1644511149
transform 1 0 47012 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_78_511
timestamp 1644511149
transform 1 0 48116 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_78_523
timestamp 1644511149
transform 1 0 49220 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_78_531
timestamp 1644511149
transform 1 0 49956 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_78_533
timestamp 1644511149
transform 1 0 50140 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_78_548
timestamp 1644511149
transform 1 0 51520 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_78_564
timestamp 1644511149
transform 1 0 52992 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_576
timestamp 1644511149
transform 1 0 54096 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_589
timestamp 1644511149
transform 1 0 55292 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_601
timestamp 1644511149
transform 1 0 56396 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_613
timestamp 1644511149
transform 1 0 57500 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_3
timestamp 1644511149
transform 1 0 1380 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_9
timestamp 1644511149
transform 1 0 1932 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_13
timestamp 1644511149
transform 1 0 2300 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_25
timestamp 1644511149
transform 1 0 3404 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_37
timestamp 1644511149
transform 1 0 4508 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_49
timestamp 1644511149
transform 1 0 5612 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_55
timestamp 1644511149
transform 1 0 6164 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_57
timestamp 1644511149
transform 1 0 6348 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_69
timestamp 1644511149
transform 1 0 7452 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_81
timestamp 1644511149
transform 1 0 8556 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_93
timestamp 1644511149
transform 1 0 9660 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_105
timestamp 1644511149
transform 1 0 10764 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_111
timestamp 1644511149
transform 1 0 11316 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_113
timestamp 1644511149
transform 1 0 11500 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_125
timestamp 1644511149
transform 1 0 12604 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_137
timestamp 1644511149
transform 1 0 13708 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_149
timestamp 1644511149
transform 1 0 14812 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_161
timestamp 1644511149
transform 1 0 15916 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_167
timestamp 1644511149
transform 1 0 16468 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_169
timestamp 1644511149
transform 1 0 16652 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_181
timestamp 1644511149
transform 1 0 17756 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_193
timestamp 1644511149
transform 1 0 18860 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_205
timestamp 1644511149
transform 1 0 19964 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_217
timestamp 1644511149
transform 1 0 21068 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_223
timestamp 1644511149
transform 1 0 21620 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_225
timestamp 1644511149
transform 1 0 21804 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_237
timestamp 1644511149
transform 1 0 22908 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_249
timestamp 1644511149
transform 1 0 24012 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_261
timestamp 1644511149
transform 1 0 25116 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_273
timestamp 1644511149
transform 1 0 26220 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_279
timestamp 1644511149
transform 1 0 26772 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_281
timestamp 1644511149
transform 1 0 26956 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_293
timestamp 1644511149
transform 1 0 28060 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_305
timestamp 1644511149
transform 1 0 29164 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_317
timestamp 1644511149
transform 1 0 30268 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_329
timestamp 1644511149
transform 1 0 31372 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_335
timestamp 1644511149
transform 1 0 31924 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_337
timestamp 1644511149
transform 1 0 32108 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_349
timestamp 1644511149
transform 1 0 33212 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_361
timestamp 1644511149
transform 1 0 34316 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_373
timestamp 1644511149
transform 1 0 35420 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_385
timestamp 1644511149
transform 1 0 36524 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_391
timestamp 1644511149
transform 1 0 37076 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_399
timestamp 1644511149
transform 1 0 37812 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_79_411
timestamp 1644511149
transform 1 0 38916 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_79_419
timestamp 1644511149
transform 1 0 39652 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_79_443
timestamp 1644511149
transform 1 0 41860 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_79_447
timestamp 1644511149
transform 1 0 42228 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_449
timestamp 1644511149
transform 1 0 42412 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_79_461
timestamp 1644511149
transform 1 0 43516 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_79_471
timestamp 1644511149
transform 1 0 44436 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_477
timestamp 1644511149
transform 1 0 44988 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_79_487
timestamp 1644511149
transform 1 0 45908 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_79_499
timestamp 1644511149
transform 1 0 47012 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_79_503
timestamp 1644511149
transform 1 0 47380 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_505
timestamp 1644511149
transform 1 0 47564 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_79_517
timestamp 1644511149
transform 1 0 48668 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_79_541
timestamp 1644511149
transform 1 0 50876 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_553
timestamp 1644511149
transform 1 0 51980 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_559
timestamp 1644511149
transform 1 0 52532 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_568
timestamp 1644511149
transform 1 0 53360 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_580
timestamp 1644511149
transform 1 0 54464 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_592
timestamp 1644511149
transform 1 0 55568 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_604
timestamp 1644511149
transform 1 0 56672 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_79_617
timestamp 1644511149
transform 1 0 57868 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_80_3
timestamp 1644511149
transform 1 0 1380 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_15
timestamp 1644511149
transform 1 0 2484 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_80_27
timestamp 1644511149
transform 1 0 3588 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_80_29
timestamp 1644511149
transform 1 0 3772 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_41
timestamp 1644511149
transform 1 0 4876 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_53
timestamp 1644511149
transform 1 0 5980 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_65
timestamp 1644511149
transform 1 0 7084 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_77
timestamp 1644511149
transform 1 0 8188 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_83
timestamp 1644511149
transform 1 0 8740 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_80_85
timestamp 1644511149
transform 1 0 8924 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_97
timestamp 1644511149
transform 1 0 10028 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_109
timestamp 1644511149
transform 1 0 11132 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_121
timestamp 1644511149
transform 1 0 12236 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_133
timestamp 1644511149
transform 1 0 13340 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_139
timestamp 1644511149
transform 1 0 13892 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_80_141
timestamp 1644511149
transform 1 0 14076 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_153
timestamp 1644511149
transform 1 0 15180 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_165
timestamp 1644511149
transform 1 0 16284 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_177
timestamp 1644511149
transform 1 0 17388 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_189
timestamp 1644511149
transform 1 0 18492 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_195
timestamp 1644511149
transform 1 0 19044 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_80_197
timestamp 1644511149
transform 1 0 19228 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_209
timestamp 1644511149
transform 1 0 20332 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_221
timestamp 1644511149
transform 1 0 21436 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_233
timestamp 1644511149
transform 1 0 22540 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_245
timestamp 1644511149
transform 1 0 23644 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_251
timestamp 1644511149
transform 1 0 24196 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_80_253
timestamp 1644511149
transform 1 0 24380 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_265
timestamp 1644511149
transform 1 0 25484 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_277
timestamp 1644511149
transform 1 0 26588 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_289
timestamp 1644511149
transform 1 0 27692 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_301
timestamp 1644511149
transform 1 0 28796 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_307
timestamp 1644511149
transform 1 0 29348 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_80_309
timestamp 1644511149
transform 1 0 29532 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_321
timestamp 1644511149
transform 1 0 30636 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_333
timestamp 1644511149
transform 1 0 31740 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_345
timestamp 1644511149
transform 1 0 32844 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_357
timestamp 1644511149
transform 1 0 33948 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_363
timestamp 1644511149
transform 1 0 34500 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_80_365
timestamp 1644511149
transform 1 0 34684 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_80_377
timestamp 1644511149
transform 1 0 35788 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_80_381
timestamp 1644511149
transform 1 0 36156 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_80_398
timestamp 1644511149
transform 1 0 37720 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_80_412
timestamp 1644511149
transform 1 0 39008 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_80_421
timestamp 1644511149
transform 1 0 39836 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_433
timestamp 1644511149
transform 1 0 40940 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_445
timestamp 1644511149
transform 1 0 42044 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_80_457
timestamp 1644511149
transform 1 0 43148 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_80_472
timestamp 1644511149
transform 1 0 44528 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_80_477
timestamp 1644511149
transform 1 0 44988 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_483
timestamp 1644511149
transform 1 0 45540 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_80_500
timestamp 1644511149
transform 1 0 47104 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_506
timestamp 1644511149
transform 1 0 47656 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_80_528
timestamp 1644511149
transform 1 0 49680 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_80_533
timestamp 1644511149
transform 1 0 50140 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_80_541
timestamp 1644511149
transform 1 0 50876 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_80_555
timestamp 1644511149
transform 1 0 52164 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_80_571
timestamp 1644511149
transform 1 0 53636 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_80_583
timestamp 1644511149
transform 1 0 54740 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_80_587
timestamp 1644511149
transform 1 0 55108 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_80_589
timestamp 1644511149
transform 1 0 55292 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_601
timestamp 1644511149
transform 1 0 56396 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_613
timestamp 1644511149
transform 1 0 57500 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_3
timestamp 1644511149
transform 1 0 1380 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_15
timestamp 1644511149
transform 1 0 2484 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_27
timestamp 1644511149
transform 1 0 3588 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_39
timestamp 1644511149
transform 1 0 4692 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_81_51
timestamp 1644511149
transform 1 0 5796 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_81_55
timestamp 1644511149
transform 1 0 6164 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_81_57
timestamp 1644511149
transform 1 0 6348 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_69
timestamp 1644511149
transform 1 0 7452 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_81
timestamp 1644511149
transform 1 0 8556 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_93
timestamp 1644511149
transform 1 0 9660 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_105
timestamp 1644511149
transform 1 0 10764 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_111
timestamp 1644511149
transform 1 0 11316 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_81_113
timestamp 1644511149
transform 1 0 11500 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_125
timestamp 1644511149
transform 1 0 12604 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_137
timestamp 1644511149
transform 1 0 13708 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_149
timestamp 1644511149
transform 1 0 14812 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_161
timestamp 1644511149
transform 1 0 15916 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_167
timestamp 1644511149
transform 1 0 16468 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_81_169
timestamp 1644511149
transform 1 0 16652 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_181
timestamp 1644511149
transform 1 0 17756 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_193
timestamp 1644511149
transform 1 0 18860 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_205
timestamp 1644511149
transform 1 0 19964 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_217
timestamp 1644511149
transform 1 0 21068 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_223
timestamp 1644511149
transform 1 0 21620 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_81_225
timestamp 1644511149
transform 1 0 21804 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_237
timestamp 1644511149
transform 1 0 22908 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_249
timestamp 1644511149
transform 1 0 24012 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_261
timestamp 1644511149
transform 1 0 25116 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_273
timestamp 1644511149
transform 1 0 26220 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_279
timestamp 1644511149
transform 1 0 26772 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_81_281
timestamp 1644511149
transform 1 0 26956 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_293
timestamp 1644511149
transform 1 0 28060 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_305
timestamp 1644511149
transform 1 0 29164 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_317
timestamp 1644511149
transform 1 0 30268 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_329
timestamp 1644511149
transform 1 0 31372 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_335
timestamp 1644511149
transform 1 0 31924 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_81_337
timestamp 1644511149
transform 1 0 32108 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_349
timestamp 1644511149
transform 1 0 33212 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_361
timestamp 1644511149
transform 1 0 34316 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_373
timestamp 1644511149
transform 1 0 35420 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_385
timestamp 1644511149
transform 1 0 36524 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_391
timestamp 1644511149
transform 1 0 37076 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_81_397
timestamp 1644511149
transform 1 0 37628 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_409
timestamp 1644511149
transform 1 0 38732 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_81_421
timestamp 1644511149
transform 1 0 39836 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_81_444
timestamp 1644511149
transform 1 0 41952 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_81_449
timestamp 1644511149
transform 1 0 42412 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_81_472
timestamp 1644511149
transform 1 0 44528 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_484
timestamp 1644511149
transform 1 0 45632 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_81_496
timestamp 1644511149
transform 1 0 46736 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_81_526
timestamp 1644511149
transform 1 0 49496 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_81_538
timestamp 1644511149
transform 1 0 50600 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_81_545
timestamp 1644511149
transform 1 0 51244 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_81_557
timestamp 1644511149
transform 1 0 52348 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_81_568
timestamp 1644511149
transform 1 0 53360 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_580
timestamp 1644511149
transform 1 0 54464 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_592
timestamp 1644511149
transform 1 0 55568 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_604
timestamp 1644511149
transform 1 0 56672 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_81_617
timestamp 1644511149
transform 1 0 57868 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_82_3
timestamp 1644511149
transform 1 0 1380 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_82_11
timestamp 1644511149
transform 1 0 2116 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_82_16
timestamp 1644511149
transform 1 0 2576 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_29
timestamp 1644511149
transform 1 0 3772 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_41
timestamp 1644511149
transform 1 0 4876 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_53
timestamp 1644511149
transform 1 0 5980 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_65
timestamp 1644511149
transform 1 0 7084 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_77
timestamp 1644511149
transform 1 0 8188 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_83
timestamp 1644511149
transform 1 0 8740 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_82_85
timestamp 1644511149
transform 1 0 8924 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_97
timestamp 1644511149
transform 1 0 10028 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_109
timestamp 1644511149
transform 1 0 11132 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_121
timestamp 1644511149
transform 1 0 12236 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_133
timestamp 1644511149
transform 1 0 13340 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_139
timestamp 1644511149
transform 1 0 13892 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_82_141
timestamp 1644511149
transform 1 0 14076 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_153
timestamp 1644511149
transform 1 0 15180 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_165
timestamp 1644511149
transform 1 0 16284 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_177
timestamp 1644511149
transform 1 0 17388 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_189
timestamp 1644511149
transform 1 0 18492 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_195
timestamp 1644511149
transform 1 0 19044 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_82_197
timestamp 1644511149
transform 1 0 19228 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_209
timestamp 1644511149
transform 1 0 20332 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_221
timestamp 1644511149
transform 1 0 21436 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_233
timestamp 1644511149
transform 1 0 22540 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_245
timestamp 1644511149
transform 1 0 23644 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_251
timestamp 1644511149
transform 1 0 24196 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_82_253
timestamp 1644511149
transform 1 0 24380 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_265
timestamp 1644511149
transform 1 0 25484 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_277
timestamp 1644511149
transform 1 0 26588 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_289
timestamp 1644511149
transform 1 0 27692 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_301
timestamp 1644511149
transform 1 0 28796 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_307
timestamp 1644511149
transform 1 0 29348 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_82_309
timestamp 1644511149
transform 1 0 29532 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_321
timestamp 1644511149
transform 1 0 30636 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_333
timestamp 1644511149
transform 1 0 31740 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_345
timestamp 1644511149
transform 1 0 32844 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_357
timestamp 1644511149
transform 1 0 33948 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_363
timestamp 1644511149
transform 1 0 34500 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_82_365
timestamp 1644511149
transform 1 0 34684 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_377
timestamp 1644511149
transform 1 0 35788 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_82_399
timestamp 1644511149
transform 1 0 37812 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_407
timestamp 1644511149
transform 1 0 38548 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_416
timestamp 1644511149
transform 1 0 39376 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_82_431
timestamp 1644511149
transform 1 0 40756 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_82_443
timestamp 1644511149
transform 1 0 41860 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_82_451
timestamp 1644511149
transform 1 0 42596 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_82_456
timestamp 1644511149
transform 1 0 43056 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_472
timestamp 1644511149
transform 1 0 44528 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_82_477
timestamp 1644511149
transform 1 0 44988 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_489
timestamp 1644511149
transform 1 0 46092 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_501
timestamp 1644511149
transform 1 0 47196 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_513
timestamp 1644511149
transform 1 0 48300 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_525
timestamp 1644511149
transform 1 0 49404 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_531
timestamp 1644511149
transform 1 0 49956 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_82_533
timestamp 1644511149
transform 1 0 50140 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_539
timestamp 1644511149
transform 1 0 50692 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_82_552
timestamp 1644511149
transform 1 0 51888 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_82_577
timestamp 1644511149
transform 1 0 54188 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_82_585
timestamp 1644511149
transform 1 0 54924 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_82_589
timestamp 1644511149
transform 1 0 55292 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_601
timestamp 1644511149
transform 1 0 56396 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_82_613
timestamp 1644511149
transform 1 0 57500 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_82_617
timestamp 1644511149
transform 1 0 57868 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_82_621
timestamp 1644511149
transform 1 0 58236 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_83_3
timestamp 1644511149
transform 1 0 1380 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_83_30
timestamp 1644511149
transform 1 0 3864 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_42
timestamp 1644511149
transform 1 0 4968 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_83_54
timestamp 1644511149
transform 1 0 6072 0 -1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_83_57
timestamp 1644511149
transform 1 0 6348 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_69
timestamp 1644511149
transform 1 0 7452 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_81
timestamp 1644511149
transform 1 0 8556 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_93
timestamp 1644511149
transform 1 0 9660 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_105
timestamp 1644511149
transform 1 0 10764 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_111
timestamp 1644511149
transform 1 0 11316 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_83_113
timestamp 1644511149
transform 1 0 11500 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_125
timestamp 1644511149
transform 1 0 12604 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_137
timestamp 1644511149
transform 1 0 13708 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_149
timestamp 1644511149
transform 1 0 14812 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_161
timestamp 1644511149
transform 1 0 15916 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_167
timestamp 1644511149
transform 1 0 16468 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_83_169
timestamp 1644511149
transform 1 0 16652 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_181
timestamp 1644511149
transform 1 0 17756 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_193
timestamp 1644511149
transform 1 0 18860 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_205
timestamp 1644511149
transform 1 0 19964 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_217
timestamp 1644511149
transform 1 0 21068 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_223
timestamp 1644511149
transform 1 0 21620 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_83_225
timestamp 1644511149
transform 1 0 21804 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_237
timestamp 1644511149
transform 1 0 22908 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_249
timestamp 1644511149
transform 1 0 24012 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_261
timestamp 1644511149
transform 1 0 25116 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_273
timestamp 1644511149
transform 1 0 26220 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_279
timestamp 1644511149
transform 1 0 26772 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_83_281
timestamp 1644511149
transform 1 0 26956 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_293
timestamp 1644511149
transform 1 0 28060 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_305
timestamp 1644511149
transform 1 0 29164 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_317
timestamp 1644511149
transform 1 0 30268 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_329
timestamp 1644511149
transform 1 0 31372 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_335
timestamp 1644511149
transform 1 0 31924 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_83_337
timestamp 1644511149
transform 1 0 32108 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_349
timestamp 1644511149
transform 1 0 33212 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_361
timestamp 1644511149
transform 1 0 34316 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_83_373
timestamp 1644511149
transform 1 0 35420 0 -1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_83_381
timestamp 1644511149
transform 1 0 36156 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_83_388
timestamp 1644511149
transform 1 0 36800 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_83_393
timestamp 1644511149
transform 1 0 37260 0 -1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_83_405
timestamp 1644511149
transform 1 0 38364 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_417
timestamp 1644511149
transform 1 0 39468 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_83_444
timestamp 1644511149
transform 1 0 41952 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_83_449
timestamp 1644511149
transform 1 0 42412 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_461
timestamp 1644511149
transform 1 0 43516 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_83_473
timestamp 1644511149
transform 1 0 44620 0 -1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_83_481
timestamp 1644511149
transform 1 0 45356 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_83_496
timestamp 1644511149
transform 1 0 46736 0 -1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_83_505
timestamp 1644511149
transform 1 0 47564 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_517
timestamp 1644511149
transform 1 0 48668 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_529
timestamp 1644511149
transform 1 0 49772 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_541
timestamp 1644511149
transform 1 0 50876 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_553
timestamp 1644511149
transform 1 0 51980 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_559
timestamp 1644511149
transform 1 0 52532 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_83_561
timestamp 1644511149
transform 1 0 52716 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_573
timestamp 1644511149
transform 1 0 53820 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_585
timestamp 1644511149
transform 1 0 54924 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_597
timestamp 1644511149
transform 1 0 56028 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_609
timestamp 1644511149
transform 1 0 57132 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_615
timestamp 1644511149
transform 1 0 57684 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_83_617
timestamp 1644511149
transform 1 0 57868 0 -1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_84_3
timestamp 1644511149
transform 1 0 1380 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_9
timestamp 1644511149
transform 1 0 1932 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_84_13
timestamp 1644511149
transform 1 0 2300 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_84_25
timestamp 1644511149
transform 1 0 3404 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_84_29
timestamp 1644511149
transform 1 0 3772 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_41
timestamp 1644511149
transform 1 0 4876 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_53
timestamp 1644511149
transform 1 0 5980 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_65
timestamp 1644511149
transform 1 0 7084 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_77
timestamp 1644511149
transform 1 0 8188 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_83
timestamp 1644511149
transform 1 0 8740 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_84_85
timestamp 1644511149
transform 1 0 8924 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_97
timestamp 1644511149
transform 1 0 10028 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_109
timestamp 1644511149
transform 1 0 11132 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_121
timestamp 1644511149
transform 1 0 12236 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_133
timestamp 1644511149
transform 1 0 13340 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_139
timestamp 1644511149
transform 1 0 13892 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_84_141
timestamp 1644511149
transform 1 0 14076 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_153
timestamp 1644511149
transform 1 0 15180 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_165
timestamp 1644511149
transform 1 0 16284 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_177
timestamp 1644511149
transform 1 0 17388 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_189
timestamp 1644511149
transform 1 0 18492 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_195
timestamp 1644511149
transform 1 0 19044 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_84_197
timestamp 1644511149
transform 1 0 19228 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_209
timestamp 1644511149
transform 1 0 20332 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_221
timestamp 1644511149
transform 1 0 21436 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_233
timestamp 1644511149
transform 1 0 22540 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_245
timestamp 1644511149
transform 1 0 23644 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_251
timestamp 1644511149
transform 1 0 24196 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_84_253
timestamp 1644511149
transform 1 0 24380 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_265
timestamp 1644511149
transform 1 0 25484 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_277
timestamp 1644511149
transform 1 0 26588 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_289
timestamp 1644511149
transform 1 0 27692 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_301
timestamp 1644511149
transform 1 0 28796 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_307
timestamp 1644511149
transform 1 0 29348 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_84_309
timestamp 1644511149
transform 1 0 29532 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_321
timestamp 1644511149
transform 1 0 30636 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_333
timestamp 1644511149
transform 1 0 31740 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_345
timestamp 1644511149
transform 1 0 32844 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_357
timestamp 1644511149
transform 1 0 33948 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_363
timestamp 1644511149
transform 1 0 34500 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_84_365
timestamp 1644511149
transform 1 0 34684 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_377
timestamp 1644511149
transform 1 0 35788 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_84_389
timestamp 1644511149
transform 1 0 36892 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_84_396
timestamp 1644511149
transform 1 0 37536 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_408
timestamp 1644511149
transform 1 0 38640 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_431
timestamp 1644511149
transform 1 0 40756 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_443
timestamp 1644511149
transform 1 0 41860 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_455
timestamp 1644511149
transform 1 0 42964 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_84_467
timestamp 1644511149
transform 1 0 44068 0 1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_84_475
timestamp 1644511149
transform 1 0 44804 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_84_477
timestamp 1644511149
transform 1 0 44988 0 1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_84_506
timestamp 1644511149
transform 1 0 47656 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_84_515
timestamp 1644511149
transform 1 0 48484 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_84_527
timestamp 1644511149
transform 1 0 49588 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_84_531
timestamp 1644511149
transform 1 0 49956 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_84_533
timestamp 1644511149
transform 1 0 50140 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_545
timestamp 1644511149
transform 1 0 51244 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_557
timestamp 1644511149
transform 1 0 52348 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_569
timestamp 1644511149
transform 1 0 53452 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_581
timestamp 1644511149
transform 1 0 54556 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_587
timestamp 1644511149
transform 1 0 55108 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_84_589
timestamp 1644511149
transform 1 0 55292 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_601
timestamp 1644511149
transform 1 0 56396 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_613
timestamp 1644511149
transform 1 0 57500 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_85_3
timestamp 1644511149
transform 1 0 1380 0 -1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_85_11
timestamp 1644511149
transform 1 0 2116 0 -1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_85_16
timestamp 1644511149
transform 1 0 2576 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_28
timestamp 1644511149
transform 1 0 3680 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_40
timestamp 1644511149
transform 1 0 4784 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_85_52
timestamp 1644511149
transform 1 0 5888 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_85_57
timestamp 1644511149
transform 1 0 6348 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_69
timestamp 1644511149
transform 1 0 7452 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_81
timestamp 1644511149
transform 1 0 8556 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_93
timestamp 1644511149
transform 1 0 9660 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_105
timestamp 1644511149
transform 1 0 10764 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_111
timestamp 1644511149
transform 1 0 11316 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_85_113
timestamp 1644511149
transform 1 0 11500 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_125
timestamp 1644511149
transform 1 0 12604 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_137
timestamp 1644511149
transform 1 0 13708 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_149
timestamp 1644511149
transform 1 0 14812 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_161
timestamp 1644511149
transform 1 0 15916 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_167
timestamp 1644511149
transform 1 0 16468 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_85_169
timestamp 1644511149
transform 1 0 16652 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_181
timestamp 1644511149
transform 1 0 17756 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_193
timestamp 1644511149
transform 1 0 18860 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_205
timestamp 1644511149
transform 1 0 19964 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_217
timestamp 1644511149
transform 1 0 21068 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_223
timestamp 1644511149
transform 1 0 21620 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_85_225
timestamp 1644511149
transform 1 0 21804 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_237
timestamp 1644511149
transform 1 0 22908 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_249
timestamp 1644511149
transform 1 0 24012 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_261
timestamp 1644511149
transform 1 0 25116 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_273
timestamp 1644511149
transform 1 0 26220 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_279
timestamp 1644511149
transform 1 0 26772 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_85_281
timestamp 1644511149
transform 1 0 26956 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_293
timestamp 1644511149
transform 1 0 28060 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_305
timestamp 1644511149
transform 1 0 29164 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_317
timestamp 1644511149
transform 1 0 30268 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_329
timestamp 1644511149
transform 1 0 31372 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_335
timestamp 1644511149
transform 1 0 31924 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_85_337
timestamp 1644511149
transform 1 0 32108 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_349
timestamp 1644511149
transform 1 0 33212 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_361
timestamp 1644511149
transform 1 0 34316 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_85_373
timestamp 1644511149
transform 1 0 35420 0 -1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_85_381
timestamp 1644511149
transform 1 0 36156 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_85_388
timestamp 1644511149
transform 1 0 36800 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_85_393
timestamp 1644511149
transform 1 0 37260 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_85_401
timestamp 1644511149
transform 1 0 37996 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_85_412
timestamp 1644511149
transform 1 0 39008 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_85_424
timestamp 1644511149
transform 1 0 40112 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_85_431
timestamp 1644511149
transform 1 0 40756 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_85_443
timestamp 1644511149
transform 1 0 41860 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_85_447
timestamp 1644511149
transform 1 0 42228 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_85_470
timestamp 1644511149
transform 1 0 44344 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_85_486
timestamp 1644511149
transform 1 0 45816 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_498
timestamp 1644511149
transform 1 0 46920 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_505
timestamp 1644511149
transform 1 0 47564 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_85_512
timestamp 1644511149
transform 1 0 48208 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_85_537
timestamp 1644511149
transform 1 0 50508 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_85_549
timestamp 1644511149
transform 1 0 51612 0 -1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_85_557
timestamp 1644511149
transform 1 0 52348 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_85_561
timestamp 1644511149
transform 1 0 52716 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_573
timestamp 1644511149
transform 1 0 53820 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_585
timestamp 1644511149
transform 1 0 54924 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_597
timestamp 1644511149
transform 1 0 56028 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_609
timestamp 1644511149
transform 1 0 57132 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_615
timestamp 1644511149
transform 1 0 57684 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_85_617
timestamp 1644511149
transform 1 0 57868 0 -1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_86_3
timestamp 1644511149
transform 1 0 1380 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_9
timestamp 1644511149
transform 1 0 1932 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_86_13
timestamp 1644511149
transform 1 0 2300 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_86_25
timestamp 1644511149
transform 1 0 3404 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_86_29
timestamp 1644511149
transform 1 0 3772 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_41
timestamp 1644511149
transform 1 0 4876 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_53
timestamp 1644511149
transform 1 0 5980 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_65
timestamp 1644511149
transform 1 0 7084 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_77
timestamp 1644511149
transform 1 0 8188 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_83
timestamp 1644511149
transform 1 0 8740 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_86_85
timestamp 1644511149
transform 1 0 8924 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_97
timestamp 1644511149
transform 1 0 10028 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_109
timestamp 1644511149
transform 1 0 11132 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_121
timestamp 1644511149
transform 1 0 12236 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_133
timestamp 1644511149
transform 1 0 13340 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_139
timestamp 1644511149
transform 1 0 13892 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_86_141
timestamp 1644511149
transform 1 0 14076 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_153
timestamp 1644511149
transform 1 0 15180 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_165
timestamp 1644511149
transform 1 0 16284 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_177
timestamp 1644511149
transform 1 0 17388 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_189
timestamp 1644511149
transform 1 0 18492 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_195
timestamp 1644511149
transform 1 0 19044 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_86_197
timestamp 1644511149
transform 1 0 19228 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_209
timestamp 1644511149
transform 1 0 20332 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_221
timestamp 1644511149
transform 1 0 21436 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_233
timestamp 1644511149
transform 1 0 22540 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_245
timestamp 1644511149
transform 1 0 23644 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_251
timestamp 1644511149
transform 1 0 24196 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_86_253
timestamp 1644511149
transform 1 0 24380 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_265
timestamp 1644511149
transform 1 0 25484 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_277
timestamp 1644511149
transform 1 0 26588 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_289
timestamp 1644511149
transform 1 0 27692 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_301
timestamp 1644511149
transform 1 0 28796 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_307
timestamp 1644511149
transform 1 0 29348 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_86_309
timestamp 1644511149
transform 1 0 29532 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_321
timestamp 1644511149
transform 1 0 30636 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_333
timestamp 1644511149
transform 1 0 31740 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_345
timestamp 1644511149
transform 1 0 32844 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_357
timestamp 1644511149
transform 1 0 33948 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_363
timestamp 1644511149
transform 1 0 34500 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_86_365
timestamp 1644511149
transform 1 0 34684 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_86_377
timestamp 1644511149
transform 1 0 35788 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_86_381
timestamp 1644511149
transform 1 0 36156 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_86_398
timestamp 1644511149
transform 1 0 37720 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_86_416
timestamp 1644511149
transform 1 0 39376 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_86_428
timestamp 1644511149
transform 1 0 40480 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_86_453
timestamp 1644511149
transform 1 0 42780 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_86_465
timestamp 1644511149
transform 1 0 43884 0 1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_86_473
timestamp 1644511149
transform 1 0 44620 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_86_498
timestamp 1644511149
transform 1 0 46920 0 1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_86_506
timestamp 1644511149
transform 1 0 47656 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_86_528
timestamp 1644511149
transform 1 0 49680 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_86_554
timestamp 1644511149
transform 1 0 52072 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_86_579
timestamp 1644511149
transform 1 0 54372 0 1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_86_587
timestamp 1644511149
transform 1 0 55108 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_86_589
timestamp 1644511149
transform 1 0 55292 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_601
timestamp 1644511149
transform 1 0 56396 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_613
timestamp 1644511149
transform 1 0 57500 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_3
timestamp 1644511149
transform 1 0 1380 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_87_30
timestamp 1644511149
transform 1 0 3864 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_42
timestamp 1644511149
transform 1 0 4968 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_87_54
timestamp 1644511149
transform 1 0 6072 0 -1 50048
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_87_57
timestamp 1644511149
transform 1 0 6348 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_69
timestamp 1644511149
transform 1 0 7452 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_81
timestamp 1644511149
transform 1 0 8556 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_93
timestamp 1644511149
transform 1 0 9660 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_105
timestamp 1644511149
transform 1 0 10764 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_111
timestamp 1644511149
transform 1 0 11316 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_87_113
timestamp 1644511149
transform 1 0 11500 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_125
timestamp 1644511149
transform 1 0 12604 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_137
timestamp 1644511149
transform 1 0 13708 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_149
timestamp 1644511149
transform 1 0 14812 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_161
timestamp 1644511149
transform 1 0 15916 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_167
timestamp 1644511149
transform 1 0 16468 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_87_169
timestamp 1644511149
transform 1 0 16652 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_181
timestamp 1644511149
transform 1 0 17756 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_193
timestamp 1644511149
transform 1 0 18860 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_205
timestamp 1644511149
transform 1 0 19964 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_217
timestamp 1644511149
transform 1 0 21068 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_223
timestamp 1644511149
transform 1 0 21620 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_87_225
timestamp 1644511149
transform 1 0 21804 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_237
timestamp 1644511149
transform 1 0 22908 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_249
timestamp 1644511149
transform 1 0 24012 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_261
timestamp 1644511149
transform 1 0 25116 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_273
timestamp 1644511149
transform 1 0 26220 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_279
timestamp 1644511149
transform 1 0 26772 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_87_281
timestamp 1644511149
transform 1 0 26956 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_293
timestamp 1644511149
transform 1 0 28060 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_305
timestamp 1644511149
transform 1 0 29164 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_317
timestamp 1644511149
transform 1 0 30268 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_329
timestamp 1644511149
transform 1 0 31372 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_335
timestamp 1644511149
transform 1 0 31924 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_87_337
timestamp 1644511149
transform 1 0 32108 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_349
timestamp 1644511149
transform 1 0 33212 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_361
timestamp 1644511149
transform 1 0 34316 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_373
timestamp 1644511149
transform 1 0 35420 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_385
timestamp 1644511149
transform 1 0 36524 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_391
timestamp 1644511149
transform 1 0 37076 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_87_393
timestamp 1644511149
transform 1 0 37260 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_399
timestamp 1644511149
transform 1 0 37812 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_87_408
timestamp 1644511149
transform 1 0 38640 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_414
timestamp 1644511149
transform 1 0 39192 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_87_420
timestamp 1644511149
transform 1 0 39744 0 -1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_87_444
timestamp 1644511149
transform 1 0 41952 0 -1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_87_449
timestamp 1644511149
transform 1 0 42412 0 -1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_87_457
timestamp 1644511149
transform 1 0 43148 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_87_479
timestamp 1644511149
transform 1 0 45172 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_491
timestamp 1644511149
transform 1 0 46276 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_87_503
timestamp 1644511149
transform 1 0 47380 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_87_521
timestamp 1644511149
transform 1 0 49036 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_87_533
timestamp 1644511149
transform 1 0 50140 0 -1 50048
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_87_556
timestamp 1644511149
transform 1 0 52256 0 -1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_87_561
timestamp 1644511149
transform 1 0 52716 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_573
timestamp 1644511149
transform 1 0 53820 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_585
timestamp 1644511149
transform 1 0 54924 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_597
timestamp 1644511149
transform 1 0 56028 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_609
timestamp 1644511149
transform 1 0 57132 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_615
timestamp 1644511149
transform 1 0 57684 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_87_617
timestamp 1644511149
transform 1 0 57868 0 -1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_88_3
timestamp 1644511149
transform 1 0 1380 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_15
timestamp 1644511149
transform 1 0 2484 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_88_27
timestamp 1644511149
transform 1 0 3588 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_88_29
timestamp 1644511149
transform 1 0 3772 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_41
timestamp 1644511149
transform 1 0 4876 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_53
timestamp 1644511149
transform 1 0 5980 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_65
timestamp 1644511149
transform 1 0 7084 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_77
timestamp 1644511149
transform 1 0 8188 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_83
timestamp 1644511149
transform 1 0 8740 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_88_85
timestamp 1644511149
transform 1 0 8924 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_97
timestamp 1644511149
transform 1 0 10028 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_109
timestamp 1644511149
transform 1 0 11132 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_121
timestamp 1644511149
transform 1 0 12236 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_133
timestamp 1644511149
transform 1 0 13340 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_139
timestamp 1644511149
transform 1 0 13892 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_88_141
timestamp 1644511149
transform 1 0 14076 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_153
timestamp 1644511149
transform 1 0 15180 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_165
timestamp 1644511149
transform 1 0 16284 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_177
timestamp 1644511149
transform 1 0 17388 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_189
timestamp 1644511149
transform 1 0 18492 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_195
timestamp 1644511149
transform 1 0 19044 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_88_197
timestamp 1644511149
transform 1 0 19228 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_209
timestamp 1644511149
transform 1 0 20332 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_221
timestamp 1644511149
transform 1 0 21436 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_233
timestamp 1644511149
transform 1 0 22540 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_245
timestamp 1644511149
transform 1 0 23644 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_251
timestamp 1644511149
transform 1 0 24196 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_88_253
timestamp 1644511149
transform 1 0 24380 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_265
timestamp 1644511149
transform 1 0 25484 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_277
timestamp 1644511149
transform 1 0 26588 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_289
timestamp 1644511149
transform 1 0 27692 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_301
timestamp 1644511149
transform 1 0 28796 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_307
timestamp 1644511149
transform 1 0 29348 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_88_309
timestamp 1644511149
transform 1 0 29532 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_321
timestamp 1644511149
transform 1 0 30636 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_333
timestamp 1644511149
transform 1 0 31740 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_345
timestamp 1644511149
transform 1 0 32844 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_357
timestamp 1644511149
transform 1 0 33948 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_363
timestamp 1644511149
transform 1 0 34500 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_88_365
timestamp 1644511149
transform 1 0 34684 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_377
timestamp 1644511149
transform 1 0 35788 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_389
timestamp 1644511149
transform 1 0 36892 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_395
timestamp 1644511149
transform 1 0 37444 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_88_412
timestamp 1644511149
transform 1 0 39008 0 1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_88_421
timestamp 1644511149
transform 1 0 39836 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_433
timestamp 1644511149
transform 1 0 40940 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_445
timestamp 1644511149
transform 1 0 42044 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_457
timestamp 1644511149
transform 1 0 43148 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_469
timestamp 1644511149
transform 1 0 44252 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_475
timestamp 1644511149
transform 1 0 44804 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_88_477
timestamp 1644511149
transform 1 0 44988 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_489
timestamp 1644511149
transform 1 0 46092 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_88_501
timestamp 1644511149
transform 1 0 47196 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_88_512
timestamp 1644511149
transform 1 0 48208 0 1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_88_522
timestamp 1644511149
transform 1 0 49128 0 1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_88_530
timestamp 1644511149
transform 1 0 49864 0 1 50048
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_88_533
timestamp 1644511149
transform 1 0 50140 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_545
timestamp 1644511149
transform 1 0 51244 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_557
timestamp 1644511149
transform 1 0 52348 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_569
timestamp 1644511149
transform 1 0 53452 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_581
timestamp 1644511149
transform 1 0 54556 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_587
timestamp 1644511149
transform 1 0 55108 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_88_589
timestamp 1644511149
transform 1 0 55292 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_601
timestamp 1644511149
transform 1 0 56396 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_613
timestamp 1644511149
transform 1 0 57500 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_3
timestamp 1644511149
transform 1 0 1380 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_15
timestamp 1644511149
transform 1 0 2484 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_27
timestamp 1644511149
transform 1 0 3588 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_39
timestamp 1644511149
transform 1 0 4692 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_89_51
timestamp 1644511149
transform 1 0 5796 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_89_55
timestamp 1644511149
transform 1 0 6164 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_89_57
timestamp 1644511149
transform 1 0 6348 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_69
timestamp 1644511149
transform 1 0 7452 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_81
timestamp 1644511149
transform 1 0 8556 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_93
timestamp 1644511149
transform 1 0 9660 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_105
timestamp 1644511149
transform 1 0 10764 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_111
timestamp 1644511149
transform 1 0 11316 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_89_113
timestamp 1644511149
transform 1 0 11500 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_125
timestamp 1644511149
transform 1 0 12604 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_137
timestamp 1644511149
transform 1 0 13708 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_149
timestamp 1644511149
transform 1 0 14812 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_161
timestamp 1644511149
transform 1 0 15916 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_167
timestamp 1644511149
transform 1 0 16468 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_89_169
timestamp 1644511149
transform 1 0 16652 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_181
timestamp 1644511149
transform 1 0 17756 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_193
timestamp 1644511149
transform 1 0 18860 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_205
timestamp 1644511149
transform 1 0 19964 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_217
timestamp 1644511149
transform 1 0 21068 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_223
timestamp 1644511149
transform 1 0 21620 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_89_225
timestamp 1644511149
transform 1 0 21804 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_237
timestamp 1644511149
transform 1 0 22908 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_249
timestamp 1644511149
transform 1 0 24012 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_261
timestamp 1644511149
transform 1 0 25116 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_273
timestamp 1644511149
transform 1 0 26220 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_279
timestamp 1644511149
transform 1 0 26772 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_89_281
timestamp 1644511149
transform 1 0 26956 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_293
timestamp 1644511149
transform 1 0 28060 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_305
timestamp 1644511149
transform 1 0 29164 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_317
timestamp 1644511149
transform 1 0 30268 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_329
timestamp 1644511149
transform 1 0 31372 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_335
timestamp 1644511149
transform 1 0 31924 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_89_337
timestamp 1644511149
transform 1 0 32108 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_349
timestamp 1644511149
transform 1 0 33212 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_361
timestamp 1644511149
transform 1 0 34316 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_373
timestamp 1644511149
transform 1 0 35420 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_385
timestamp 1644511149
transform 1 0 36524 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_391
timestamp 1644511149
transform 1 0 37076 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_89_393
timestamp 1644511149
transform 1 0 37260 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_405
timestamp 1644511149
transform 1 0 38364 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_417
timestamp 1644511149
transform 1 0 39468 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_429
timestamp 1644511149
transform 1 0 40572 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_441
timestamp 1644511149
transform 1 0 41676 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_447
timestamp 1644511149
transform 1 0 42228 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_89_449
timestamp 1644511149
transform 1 0 42412 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_461
timestamp 1644511149
transform 1 0 43516 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_89_473
timestamp 1644511149
transform 1 0 44620 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_89_477
timestamp 1644511149
transform 1 0 44988 0 -1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_89_485
timestamp 1644511149
transform 1 0 45724 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_89_489
timestamp 1644511149
transform 1 0 46092 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_89_501
timestamp 1644511149
transform 1 0 47196 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_89_505
timestamp 1644511149
transform 1 0 47564 0 -1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_89_513
timestamp 1644511149
transform 1 0 48300 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_89_517
timestamp 1644511149
transform 1 0 48668 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_89_526
timestamp 1644511149
transform 1 0 49496 0 -1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_89_537
timestamp 1644511149
transform 1 0 50508 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_89_549
timestamp 1644511149
transform 1 0 51612 0 -1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_89_557
timestamp 1644511149
transform 1 0 52348 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_89_561
timestamp 1644511149
transform 1 0 52716 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_573
timestamp 1644511149
transform 1 0 53820 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_585
timestamp 1644511149
transform 1 0 54924 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_597
timestamp 1644511149
transform 1 0 56028 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_609
timestamp 1644511149
transform 1 0 57132 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_615
timestamp 1644511149
transform 1 0 57684 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_89_617
timestamp 1644511149
transform 1 0 57868 0 -1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_90_3
timestamp 1644511149
transform 1 0 1380 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_15
timestamp 1644511149
transform 1 0 2484 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_90_27
timestamp 1644511149
transform 1 0 3588 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_90_29
timestamp 1644511149
transform 1 0 3772 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_41
timestamp 1644511149
transform 1 0 4876 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_53
timestamp 1644511149
transform 1 0 5980 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_65
timestamp 1644511149
transform 1 0 7084 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_77
timestamp 1644511149
transform 1 0 8188 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_83
timestamp 1644511149
transform 1 0 8740 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_90_85
timestamp 1644511149
transform 1 0 8924 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_97
timestamp 1644511149
transform 1 0 10028 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_109
timestamp 1644511149
transform 1 0 11132 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_121
timestamp 1644511149
transform 1 0 12236 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_133
timestamp 1644511149
transform 1 0 13340 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_139
timestamp 1644511149
transform 1 0 13892 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_90_141
timestamp 1644511149
transform 1 0 14076 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_153
timestamp 1644511149
transform 1 0 15180 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_165
timestamp 1644511149
transform 1 0 16284 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_177
timestamp 1644511149
transform 1 0 17388 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_189
timestamp 1644511149
transform 1 0 18492 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_195
timestamp 1644511149
transform 1 0 19044 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_90_197
timestamp 1644511149
transform 1 0 19228 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_209
timestamp 1644511149
transform 1 0 20332 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_221
timestamp 1644511149
transform 1 0 21436 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_233
timestamp 1644511149
transform 1 0 22540 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_245
timestamp 1644511149
transform 1 0 23644 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_251
timestamp 1644511149
transform 1 0 24196 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_90_253
timestamp 1644511149
transform 1 0 24380 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_265
timestamp 1644511149
transform 1 0 25484 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_277
timestamp 1644511149
transform 1 0 26588 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_289
timestamp 1644511149
transform 1 0 27692 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_301
timestamp 1644511149
transform 1 0 28796 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_307
timestamp 1644511149
transform 1 0 29348 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_90_309
timestamp 1644511149
transform 1 0 29532 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_321
timestamp 1644511149
transform 1 0 30636 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_333
timestamp 1644511149
transform 1 0 31740 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_345
timestamp 1644511149
transform 1 0 32844 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_357
timestamp 1644511149
transform 1 0 33948 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_363
timestamp 1644511149
transform 1 0 34500 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_90_365
timestamp 1644511149
transform 1 0 34684 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_377
timestamp 1644511149
transform 1 0 35788 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_389
timestamp 1644511149
transform 1 0 36892 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_401
timestamp 1644511149
transform 1 0 37996 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_413
timestamp 1644511149
transform 1 0 39100 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_419
timestamp 1644511149
transform 1 0 39652 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_90_421
timestamp 1644511149
transform 1 0 39836 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_433
timestamp 1644511149
transform 1 0 40940 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_445
timestamp 1644511149
transform 1 0 42044 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_457
timestamp 1644511149
transform 1 0 43148 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_469
timestamp 1644511149
transform 1 0 44252 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_475
timestamp 1644511149
transform 1 0 44804 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_90_480
timestamp 1644511149
transform 1 0 45264 0 1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_90_493
timestamp 1644511149
transform 1 0 46460 0 1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_90_501
timestamp 1644511149
transform 1 0 47196 0 1 51136
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_90_508
timestamp 1644511149
transform 1 0 47840 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_520
timestamp 1644511149
transform 1 0 48944 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_90_533
timestamp 1644511149
transform 1 0 50140 0 1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_90_537
timestamp 1644511149
transform 1 0 50508 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_90_541
timestamp 1644511149
transform 1 0 50876 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_553
timestamp 1644511149
transform 1 0 51980 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_565
timestamp 1644511149
transform 1 0 53084 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_90_577
timestamp 1644511149
transform 1 0 54188 0 1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_90_585
timestamp 1644511149
transform 1 0 54924 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_90_589
timestamp 1644511149
transform 1 0 55292 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_601
timestamp 1644511149
transform 1 0 56396 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_613
timestamp 1644511149
transform 1 0 57500 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_3
timestamp 1644511149
transform 1 0 1380 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_15
timestamp 1644511149
transform 1 0 2484 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_27
timestamp 1644511149
transform 1 0 3588 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_39
timestamp 1644511149
transform 1 0 4692 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_91_51
timestamp 1644511149
transform 1 0 5796 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_91_55
timestamp 1644511149
transform 1 0 6164 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_91_57
timestamp 1644511149
transform 1 0 6348 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_69
timestamp 1644511149
transform 1 0 7452 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_81
timestamp 1644511149
transform 1 0 8556 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_93
timestamp 1644511149
transform 1 0 9660 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_105
timestamp 1644511149
transform 1 0 10764 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_111
timestamp 1644511149
transform 1 0 11316 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_91_113
timestamp 1644511149
transform 1 0 11500 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_125
timestamp 1644511149
transform 1 0 12604 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_137
timestamp 1644511149
transform 1 0 13708 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_149
timestamp 1644511149
transform 1 0 14812 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_161
timestamp 1644511149
transform 1 0 15916 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_167
timestamp 1644511149
transform 1 0 16468 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_91_169
timestamp 1644511149
transform 1 0 16652 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_181
timestamp 1644511149
transform 1 0 17756 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_193
timestamp 1644511149
transform 1 0 18860 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_205
timestamp 1644511149
transform 1 0 19964 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_217
timestamp 1644511149
transform 1 0 21068 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_223
timestamp 1644511149
transform 1 0 21620 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_91_225
timestamp 1644511149
transform 1 0 21804 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_237
timestamp 1644511149
transform 1 0 22908 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_249
timestamp 1644511149
transform 1 0 24012 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_261
timestamp 1644511149
transform 1 0 25116 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_273
timestamp 1644511149
transform 1 0 26220 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_279
timestamp 1644511149
transform 1 0 26772 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_91_281
timestamp 1644511149
transform 1 0 26956 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_293
timestamp 1644511149
transform 1 0 28060 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_305
timestamp 1644511149
transform 1 0 29164 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_317
timestamp 1644511149
transform 1 0 30268 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_329
timestamp 1644511149
transform 1 0 31372 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_335
timestamp 1644511149
transform 1 0 31924 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_91_337
timestamp 1644511149
transform 1 0 32108 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_349
timestamp 1644511149
transform 1 0 33212 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_361
timestamp 1644511149
transform 1 0 34316 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_373
timestamp 1644511149
transform 1 0 35420 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_385
timestamp 1644511149
transform 1 0 36524 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_391
timestamp 1644511149
transform 1 0 37076 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_91_393
timestamp 1644511149
transform 1 0 37260 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_405
timestamp 1644511149
transform 1 0 38364 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_417
timestamp 1644511149
transform 1 0 39468 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_429
timestamp 1644511149
transform 1 0 40572 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_441
timestamp 1644511149
transform 1 0 41676 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_447
timestamp 1644511149
transform 1 0 42228 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_91_470
timestamp 1644511149
transform 1 0 44344 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_91_482
timestamp 1644511149
transform 1 0 45448 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_91_489
timestamp 1644511149
transform 1 0 46092 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_91_499
timestamp 1644511149
transform 1 0 47012 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_91_503
timestamp 1644511149
transform 1 0 47380 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_91_510
timestamp 1644511149
transform 1 0 48024 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_91_522
timestamp 1644511149
transform 1 0 49128 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_91_533
timestamp 1644511149
transform 1 0 50140 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_91_544
timestamp 1644511149
transform 1 0 51152 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_91_551
timestamp 1644511149
transform 1 0 51796 0 -1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_91_559
timestamp 1644511149
transform 1 0 52532 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_91_561
timestamp 1644511149
transform 1 0 52716 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_573
timestamp 1644511149
transform 1 0 53820 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_585
timestamp 1644511149
transform 1 0 54924 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_597
timestamp 1644511149
transform 1 0 56028 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_609
timestamp 1644511149
transform 1 0 57132 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_615
timestamp 1644511149
transform 1 0 57684 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_91_617
timestamp 1644511149
transform 1 0 57868 0 -1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_92_3
timestamp 1644511149
transform 1 0 1380 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_15
timestamp 1644511149
transform 1 0 2484 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_92_27
timestamp 1644511149
transform 1 0 3588 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_92_29
timestamp 1644511149
transform 1 0 3772 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_41
timestamp 1644511149
transform 1 0 4876 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_53
timestamp 1644511149
transform 1 0 5980 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_65
timestamp 1644511149
transform 1 0 7084 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_77
timestamp 1644511149
transform 1 0 8188 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_83
timestamp 1644511149
transform 1 0 8740 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_92_85
timestamp 1644511149
transform 1 0 8924 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_97
timestamp 1644511149
transform 1 0 10028 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_109
timestamp 1644511149
transform 1 0 11132 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_121
timestamp 1644511149
transform 1 0 12236 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_133
timestamp 1644511149
transform 1 0 13340 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_139
timestamp 1644511149
transform 1 0 13892 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_92_141
timestamp 1644511149
transform 1 0 14076 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_153
timestamp 1644511149
transform 1 0 15180 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_165
timestamp 1644511149
transform 1 0 16284 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_177
timestamp 1644511149
transform 1 0 17388 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_189
timestamp 1644511149
transform 1 0 18492 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_195
timestamp 1644511149
transform 1 0 19044 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_92_197
timestamp 1644511149
transform 1 0 19228 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_209
timestamp 1644511149
transform 1 0 20332 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_221
timestamp 1644511149
transform 1 0 21436 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_233
timestamp 1644511149
transform 1 0 22540 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_245
timestamp 1644511149
transform 1 0 23644 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_251
timestamp 1644511149
transform 1 0 24196 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_92_253
timestamp 1644511149
transform 1 0 24380 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_265
timestamp 1644511149
transform 1 0 25484 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_277
timestamp 1644511149
transform 1 0 26588 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_289
timestamp 1644511149
transform 1 0 27692 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_301
timestamp 1644511149
transform 1 0 28796 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_307
timestamp 1644511149
transform 1 0 29348 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_92_309
timestamp 1644511149
transform 1 0 29532 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_321
timestamp 1644511149
transform 1 0 30636 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_333
timestamp 1644511149
transform 1 0 31740 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_345
timestamp 1644511149
transform 1 0 32844 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_357
timestamp 1644511149
transform 1 0 33948 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_363
timestamp 1644511149
transform 1 0 34500 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_92_365
timestamp 1644511149
transform 1 0 34684 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_377
timestamp 1644511149
transform 1 0 35788 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_389
timestamp 1644511149
transform 1 0 36892 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_401
timestamp 1644511149
transform 1 0 37996 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_413
timestamp 1644511149
transform 1 0 39100 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_419
timestamp 1644511149
transform 1 0 39652 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_92_421
timestamp 1644511149
transform 1 0 39836 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_92_433
timestamp 1644511149
transform 1 0 40940 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_92_439
timestamp 1644511149
transform 1 0 41492 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_92_464
timestamp 1644511149
transform 1 0 43792 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_92_471
timestamp 1644511149
transform 1 0 44436 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_92_475
timestamp 1644511149
transform 1 0 44804 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_92_493
timestamp 1644511149
transform 1 0 46460 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_92_500
timestamp 1644511149
transform 1 0 47104 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_92_520
timestamp 1644511149
transform 1 0 48944 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_92_528
timestamp 1644511149
transform 1 0 49680 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_92_543
timestamp 1644511149
transform 1 0 51060 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_555
timestamp 1644511149
transform 1 0 52164 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_567
timestamp 1644511149
transform 1 0 53268 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_92_579
timestamp 1644511149
transform 1 0 54372 0 1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_92_587
timestamp 1644511149
transform 1 0 55108 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_92_589
timestamp 1644511149
transform 1 0 55292 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_601
timestamp 1644511149
transform 1 0 56396 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_613
timestamp 1644511149
transform 1 0 57500 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_3
timestamp 1644511149
transform 1 0 1380 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_15
timestamp 1644511149
transform 1 0 2484 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_27
timestamp 1644511149
transform 1 0 3588 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_39
timestamp 1644511149
transform 1 0 4692 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_93_51
timestamp 1644511149
transform 1 0 5796 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_93_55
timestamp 1644511149
transform 1 0 6164 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_93_57
timestamp 1644511149
transform 1 0 6348 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_69
timestamp 1644511149
transform 1 0 7452 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_81
timestamp 1644511149
transform 1 0 8556 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_93
timestamp 1644511149
transform 1 0 9660 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_105
timestamp 1644511149
transform 1 0 10764 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_111
timestamp 1644511149
transform 1 0 11316 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_93_113
timestamp 1644511149
transform 1 0 11500 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_125
timestamp 1644511149
transform 1 0 12604 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_137
timestamp 1644511149
transform 1 0 13708 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_149
timestamp 1644511149
transform 1 0 14812 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_161
timestamp 1644511149
transform 1 0 15916 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_167
timestamp 1644511149
transform 1 0 16468 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_93_169
timestamp 1644511149
transform 1 0 16652 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_181
timestamp 1644511149
transform 1 0 17756 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_193
timestamp 1644511149
transform 1 0 18860 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_205
timestamp 1644511149
transform 1 0 19964 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_217
timestamp 1644511149
transform 1 0 21068 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_223
timestamp 1644511149
transform 1 0 21620 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_93_225
timestamp 1644511149
transform 1 0 21804 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_237
timestamp 1644511149
transform 1 0 22908 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_249
timestamp 1644511149
transform 1 0 24012 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_261
timestamp 1644511149
transform 1 0 25116 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_273
timestamp 1644511149
transform 1 0 26220 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_279
timestamp 1644511149
transform 1 0 26772 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_93_281
timestamp 1644511149
transform 1 0 26956 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_293
timestamp 1644511149
transform 1 0 28060 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_305
timestamp 1644511149
transform 1 0 29164 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_317
timestamp 1644511149
transform 1 0 30268 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_329
timestamp 1644511149
transform 1 0 31372 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_335
timestamp 1644511149
transform 1 0 31924 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_93_337
timestamp 1644511149
transform 1 0 32108 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_349
timestamp 1644511149
transform 1 0 33212 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_361
timestamp 1644511149
transform 1 0 34316 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_373
timestamp 1644511149
transform 1 0 35420 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_385
timestamp 1644511149
transform 1 0 36524 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_391
timestamp 1644511149
transform 1 0 37076 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_93_393
timestamp 1644511149
transform 1 0 37260 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_405
timestamp 1644511149
transform 1 0 38364 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_417
timestamp 1644511149
transform 1 0 39468 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_429
timestamp 1644511149
transform 1 0 40572 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_441
timestamp 1644511149
transform 1 0 41676 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_447
timestamp 1644511149
transform 1 0 42228 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_93_470
timestamp 1644511149
transform 1 0 44344 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_498
timestamp 1644511149
transform 1 0 46920 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_93_505
timestamp 1644511149
transform 1 0 47564 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_93_511
timestamp 1644511149
transform 1 0 48116 0 -1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_93_519
timestamp 1644511149
transform 1 0 48852 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_93_524
timestamp 1644511149
transform 1 0 49312 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_93_538
timestamp 1644511149
transform 1 0 50600 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_93_550
timestamp 1644511149
transform 1 0 51704 0 -1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_93_558
timestamp 1644511149
transform 1 0 52440 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_93_561
timestamp 1644511149
transform 1 0 52716 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_573
timestamp 1644511149
transform 1 0 53820 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_585
timestamp 1644511149
transform 1 0 54924 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_597
timestamp 1644511149
transform 1 0 56028 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_609
timestamp 1644511149
transform 1 0 57132 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_615
timestamp 1644511149
transform 1 0 57684 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_93_617
timestamp 1644511149
transform 1 0 57868 0 -1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_94_3
timestamp 1644511149
transform 1 0 1380 0 1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_94_11
timestamp 1644511149
transform 1 0 2116 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_94_16
timestamp 1644511149
transform 1 0 2576 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_29
timestamp 1644511149
transform 1 0 3772 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_41
timestamp 1644511149
transform 1 0 4876 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_53
timestamp 1644511149
transform 1 0 5980 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_65
timestamp 1644511149
transform 1 0 7084 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_77
timestamp 1644511149
transform 1 0 8188 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_83
timestamp 1644511149
transform 1 0 8740 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_94_85
timestamp 1644511149
transform 1 0 8924 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_97
timestamp 1644511149
transform 1 0 10028 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_109
timestamp 1644511149
transform 1 0 11132 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_121
timestamp 1644511149
transform 1 0 12236 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_133
timestamp 1644511149
transform 1 0 13340 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_139
timestamp 1644511149
transform 1 0 13892 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_94_141
timestamp 1644511149
transform 1 0 14076 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_153
timestamp 1644511149
transform 1 0 15180 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_165
timestamp 1644511149
transform 1 0 16284 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_177
timestamp 1644511149
transform 1 0 17388 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_189
timestamp 1644511149
transform 1 0 18492 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_195
timestamp 1644511149
transform 1 0 19044 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_94_197
timestamp 1644511149
transform 1 0 19228 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_209
timestamp 1644511149
transform 1 0 20332 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_221
timestamp 1644511149
transform 1 0 21436 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_233
timestamp 1644511149
transform 1 0 22540 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_245
timestamp 1644511149
transform 1 0 23644 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_251
timestamp 1644511149
transform 1 0 24196 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_94_253
timestamp 1644511149
transform 1 0 24380 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_265
timestamp 1644511149
transform 1 0 25484 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_277
timestamp 1644511149
transform 1 0 26588 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_289
timestamp 1644511149
transform 1 0 27692 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_301
timestamp 1644511149
transform 1 0 28796 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_307
timestamp 1644511149
transform 1 0 29348 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_94_309
timestamp 1644511149
transform 1 0 29532 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_321
timestamp 1644511149
transform 1 0 30636 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_333
timestamp 1644511149
transform 1 0 31740 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_345
timestamp 1644511149
transform 1 0 32844 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_357
timestamp 1644511149
transform 1 0 33948 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_363
timestamp 1644511149
transform 1 0 34500 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_94_365
timestamp 1644511149
transform 1 0 34684 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_377
timestamp 1644511149
transform 1 0 35788 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_389
timestamp 1644511149
transform 1 0 36892 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_401
timestamp 1644511149
transform 1 0 37996 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_413
timestamp 1644511149
transform 1 0 39100 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_419
timestamp 1644511149
transform 1 0 39652 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_94_421
timestamp 1644511149
transform 1 0 39836 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_433
timestamp 1644511149
transform 1 0 40940 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_94_445
timestamp 1644511149
transform 1 0 42044 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_94_452
timestamp 1644511149
transform 1 0 42688 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_464
timestamp 1644511149
transform 1 0 43792 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_94_477
timestamp 1644511149
transform 1 0 44988 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_94_481
timestamp 1644511149
transform 1 0 45356 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_94_486
timestamp 1644511149
transform 1 0 45816 0 1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_94_497
timestamp 1644511149
transform 1 0 46828 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_509
timestamp 1644511149
transform 1 0 47932 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_94_521
timestamp 1644511149
transform 1 0 49036 0 1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_94_529
timestamp 1644511149
transform 1 0 49772 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_94_533
timestamp 1644511149
transform 1 0 50140 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_545
timestamp 1644511149
transform 1 0 51244 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_557
timestamp 1644511149
transform 1 0 52348 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_569
timestamp 1644511149
transform 1 0 53452 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_581
timestamp 1644511149
transform 1 0 54556 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_587
timestamp 1644511149
transform 1 0 55108 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_94_589
timestamp 1644511149
transform 1 0 55292 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_601
timestamp 1644511149
transform 1 0 56396 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_613
timestamp 1644511149
transform 1 0 57500 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_3
timestamp 1644511149
transform 1 0 1380 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_95_30
timestamp 1644511149
transform 1 0 3864 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_42
timestamp 1644511149
transform 1 0 4968 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_95_54
timestamp 1644511149
transform 1 0 6072 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_95_57
timestamp 1644511149
transform 1 0 6348 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_69
timestamp 1644511149
transform 1 0 7452 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_81
timestamp 1644511149
transform 1 0 8556 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_93
timestamp 1644511149
transform 1 0 9660 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_105
timestamp 1644511149
transform 1 0 10764 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_111
timestamp 1644511149
transform 1 0 11316 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_95_113
timestamp 1644511149
transform 1 0 11500 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_125
timestamp 1644511149
transform 1 0 12604 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_137
timestamp 1644511149
transform 1 0 13708 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_149
timestamp 1644511149
transform 1 0 14812 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_161
timestamp 1644511149
transform 1 0 15916 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_167
timestamp 1644511149
transform 1 0 16468 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_95_169
timestamp 1644511149
transform 1 0 16652 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_181
timestamp 1644511149
transform 1 0 17756 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_193
timestamp 1644511149
transform 1 0 18860 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_205
timestamp 1644511149
transform 1 0 19964 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_217
timestamp 1644511149
transform 1 0 21068 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_223
timestamp 1644511149
transform 1 0 21620 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_95_225
timestamp 1644511149
transform 1 0 21804 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_237
timestamp 1644511149
transform 1 0 22908 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_249
timestamp 1644511149
transform 1 0 24012 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_261
timestamp 1644511149
transform 1 0 25116 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_273
timestamp 1644511149
transform 1 0 26220 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_279
timestamp 1644511149
transform 1 0 26772 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_95_281
timestamp 1644511149
transform 1 0 26956 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_293
timestamp 1644511149
transform 1 0 28060 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_305
timestamp 1644511149
transform 1 0 29164 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_317
timestamp 1644511149
transform 1 0 30268 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_329
timestamp 1644511149
transform 1 0 31372 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_335
timestamp 1644511149
transform 1 0 31924 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_95_337
timestamp 1644511149
transform 1 0 32108 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_349
timestamp 1644511149
transform 1 0 33212 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_361
timestamp 1644511149
transform 1 0 34316 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_373
timestamp 1644511149
transform 1 0 35420 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_385
timestamp 1644511149
transform 1 0 36524 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_391
timestamp 1644511149
transform 1 0 37076 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_95_393
timestamp 1644511149
transform 1 0 37260 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_405
timestamp 1644511149
transform 1 0 38364 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_417
timestamp 1644511149
transform 1 0 39468 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_429
timestamp 1644511149
transform 1 0 40572 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_441
timestamp 1644511149
transform 1 0 41676 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_447
timestamp 1644511149
transform 1 0 42228 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_95_449
timestamp 1644511149
transform 1 0 42412 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_461
timestamp 1644511149
transform 1 0 43516 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_473
timestamp 1644511149
transform 1 0 44620 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_485
timestamp 1644511149
transform 1 0 45724 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_95_494
timestamp 1644511149
transform 1 0 46552 0 -1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_95_502
timestamp 1644511149
transform 1 0 47288 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_95_505
timestamp 1644511149
transform 1 0 47564 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_517
timestamp 1644511149
transform 1 0 48668 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_529
timestamp 1644511149
transform 1 0 49772 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_541
timestamp 1644511149
transform 1 0 50876 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_553
timestamp 1644511149
transform 1 0 51980 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_559
timestamp 1644511149
transform 1 0 52532 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_95_561
timestamp 1644511149
transform 1 0 52716 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_573
timestamp 1644511149
transform 1 0 53820 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_585
timestamp 1644511149
transform 1 0 54924 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_597
timestamp 1644511149
transform 1 0 56028 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_609
timestamp 1644511149
transform 1 0 57132 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_615
timestamp 1644511149
transform 1 0 57684 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_95_617
timestamp 1644511149
transform 1 0 57868 0 -1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_96_3
timestamp 1644511149
transform 1 0 1380 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_9
timestamp 1644511149
transform 1 0 1932 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_96_13
timestamp 1644511149
transform 1 0 2300 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_96_25
timestamp 1644511149
transform 1 0 3404 0 1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_96_29
timestamp 1644511149
transform 1 0 3772 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_41
timestamp 1644511149
transform 1 0 4876 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_53
timestamp 1644511149
transform 1 0 5980 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_65
timestamp 1644511149
transform 1 0 7084 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_77
timestamp 1644511149
transform 1 0 8188 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_83
timestamp 1644511149
transform 1 0 8740 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_96_85
timestamp 1644511149
transform 1 0 8924 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_97
timestamp 1644511149
transform 1 0 10028 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_109
timestamp 1644511149
transform 1 0 11132 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_121
timestamp 1644511149
transform 1 0 12236 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_133
timestamp 1644511149
transform 1 0 13340 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_139
timestamp 1644511149
transform 1 0 13892 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_96_141
timestamp 1644511149
transform 1 0 14076 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_153
timestamp 1644511149
transform 1 0 15180 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_165
timestamp 1644511149
transform 1 0 16284 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_177
timestamp 1644511149
transform 1 0 17388 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_189
timestamp 1644511149
transform 1 0 18492 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_195
timestamp 1644511149
transform 1 0 19044 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_96_197
timestamp 1644511149
transform 1 0 19228 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_209
timestamp 1644511149
transform 1 0 20332 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_221
timestamp 1644511149
transform 1 0 21436 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_233
timestamp 1644511149
transform 1 0 22540 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_245
timestamp 1644511149
transform 1 0 23644 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_251
timestamp 1644511149
transform 1 0 24196 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_96_253
timestamp 1644511149
transform 1 0 24380 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_265
timestamp 1644511149
transform 1 0 25484 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_277
timestamp 1644511149
transform 1 0 26588 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_289
timestamp 1644511149
transform 1 0 27692 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_301
timestamp 1644511149
transform 1 0 28796 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_307
timestamp 1644511149
transform 1 0 29348 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_96_309
timestamp 1644511149
transform 1 0 29532 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_321
timestamp 1644511149
transform 1 0 30636 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_333
timestamp 1644511149
transform 1 0 31740 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_345
timestamp 1644511149
transform 1 0 32844 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_357
timestamp 1644511149
transform 1 0 33948 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_363
timestamp 1644511149
transform 1 0 34500 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_96_365
timestamp 1644511149
transform 1 0 34684 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_377
timestamp 1644511149
transform 1 0 35788 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_389
timestamp 1644511149
transform 1 0 36892 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_401
timestamp 1644511149
transform 1 0 37996 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_413
timestamp 1644511149
transform 1 0 39100 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_419
timestamp 1644511149
transform 1 0 39652 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_96_421
timestamp 1644511149
transform 1 0 39836 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_433
timestamp 1644511149
transform 1 0 40940 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_96_445
timestamp 1644511149
transform 1 0 42044 0 1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_96_469
timestamp 1644511149
transform 1 0 44252 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_475
timestamp 1644511149
transform 1 0 44804 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_96_477
timestamp 1644511149
transform 1 0 44988 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_489
timestamp 1644511149
transform 1 0 46092 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_501
timestamp 1644511149
transform 1 0 47196 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_513
timestamp 1644511149
transform 1 0 48300 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_525
timestamp 1644511149
transform 1 0 49404 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_531
timestamp 1644511149
transform 1 0 49956 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_96_533
timestamp 1644511149
transform 1 0 50140 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_545
timestamp 1644511149
transform 1 0 51244 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_557
timestamp 1644511149
transform 1 0 52348 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_569
timestamp 1644511149
transform 1 0 53452 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_581
timestamp 1644511149
transform 1 0 54556 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_587
timestamp 1644511149
transform 1 0 55108 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_96_589
timestamp 1644511149
transform 1 0 55292 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_601
timestamp 1644511149
transform 1 0 56396 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_613
timestamp 1644511149
transform 1 0 57500 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_3
timestamp 1644511149
transform 1 0 1380 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_15
timestamp 1644511149
transform 1 0 2484 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_27
timestamp 1644511149
transform 1 0 3588 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_39
timestamp 1644511149
transform 1 0 4692 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_97_51
timestamp 1644511149
transform 1 0 5796 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_97_55
timestamp 1644511149
transform 1 0 6164 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_97_57
timestamp 1644511149
transform 1 0 6348 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_69
timestamp 1644511149
transform 1 0 7452 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_97_81
timestamp 1644511149
transform 1 0 8556 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_97_85
timestamp 1644511149
transform 1 0 8924 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_97_89
timestamp 1644511149
transform 1 0 9292 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_97_101
timestamp 1644511149
transform 1 0 10396 0 -1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_97_109
timestamp 1644511149
transform 1 0 11132 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_97_113
timestamp 1644511149
transform 1 0 11500 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_125
timestamp 1644511149
transform 1 0 12604 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_137
timestamp 1644511149
transform 1 0 13708 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_149
timestamp 1644511149
transform 1 0 14812 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_161
timestamp 1644511149
transform 1 0 15916 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_167
timestamp 1644511149
transform 1 0 16468 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_97_169
timestamp 1644511149
transform 1 0 16652 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_181
timestamp 1644511149
transform 1 0 17756 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_193
timestamp 1644511149
transform 1 0 18860 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_205
timestamp 1644511149
transform 1 0 19964 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_217
timestamp 1644511149
transform 1 0 21068 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_223
timestamp 1644511149
transform 1 0 21620 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_97_225
timestamp 1644511149
transform 1 0 21804 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_237
timestamp 1644511149
transform 1 0 22908 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_249
timestamp 1644511149
transform 1 0 24012 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_97_261
timestamp 1644511149
transform 1 0 25116 0 -1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_97_269
timestamp 1644511149
transform 1 0 25852 0 -1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_97_274
timestamp 1644511149
transform 1 0 26312 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_97_281
timestamp 1644511149
transform 1 0 26956 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_293
timestamp 1644511149
transform 1 0 28060 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_305
timestamp 1644511149
transform 1 0 29164 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_317
timestamp 1644511149
transform 1 0 30268 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_329
timestamp 1644511149
transform 1 0 31372 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_335
timestamp 1644511149
transform 1 0 31924 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_97_337
timestamp 1644511149
transform 1 0 32108 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_349
timestamp 1644511149
transform 1 0 33212 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_361
timestamp 1644511149
transform 1 0 34316 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_97_373
timestamp 1644511149
transform 1 0 35420 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_97_380
timestamp 1644511149
transform 1 0 36064 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_393
timestamp 1644511149
transform 1 0 37260 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_405
timestamp 1644511149
transform 1 0 38364 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_417
timestamp 1644511149
transform 1 0 39468 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_429
timestamp 1644511149
transform 1 0 40572 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_441
timestamp 1644511149
transform 1 0 41676 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_447
timestamp 1644511149
transform 1 0 42228 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_97_470
timestamp 1644511149
transform 1 0 44344 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_482
timestamp 1644511149
transform 1 0 45448 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_97_494
timestamp 1644511149
transform 1 0 46552 0 -1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_97_502
timestamp 1644511149
transform 1 0 47288 0 -1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_97_505
timestamp 1644511149
transform 1 0 47564 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_517
timestamp 1644511149
transform 1 0 48668 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_529
timestamp 1644511149
transform 1 0 49772 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_541
timestamp 1644511149
transform 1 0 50876 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_553
timestamp 1644511149
transform 1 0 51980 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_559
timestamp 1644511149
transform 1 0 52532 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_97_561
timestamp 1644511149
transform 1 0 52716 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_573
timestamp 1644511149
transform 1 0 53820 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_585
timestamp 1644511149
transform 1 0 54924 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_597
timestamp 1644511149
transform 1 0 56028 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_609
timestamp 1644511149
transform 1 0 57132 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_615
timestamp 1644511149
transform 1 0 57684 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_97_617
timestamp 1644511149
transform 1 0 57868 0 -1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_98_3
timestamp 1644511149
transform 1 0 1380 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_15
timestamp 1644511149
transform 1 0 2484 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_98_27
timestamp 1644511149
transform 1 0 3588 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_98_29
timestamp 1644511149
transform 1 0 3772 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_41
timestamp 1644511149
transform 1 0 4876 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_53
timestamp 1644511149
transform 1 0 5980 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_65
timestamp 1644511149
transform 1 0 7084 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_77
timestamp 1644511149
transform 1 0 8188 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_83
timestamp 1644511149
transform 1 0 8740 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_98_85
timestamp 1644511149
transform 1 0 8924 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_97
timestamp 1644511149
transform 1 0 10028 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_109
timestamp 1644511149
transform 1 0 11132 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_121
timestamp 1644511149
transform 1 0 12236 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_133
timestamp 1644511149
transform 1 0 13340 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_139
timestamp 1644511149
transform 1 0 13892 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_98_141
timestamp 1644511149
transform 1 0 14076 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_153
timestamp 1644511149
transform 1 0 15180 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_165
timestamp 1644511149
transform 1 0 16284 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_177
timestamp 1644511149
transform 1 0 17388 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_189
timestamp 1644511149
transform 1 0 18492 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_195
timestamp 1644511149
transform 1 0 19044 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_98_197
timestamp 1644511149
transform 1 0 19228 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_209
timestamp 1644511149
transform 1 0 20332 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_221
timestamp 1644511149
transform 1 0 21436 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_233
timestamp 1644511149
transform 1 0 22540 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_245
timestamp 1644511149
transform 1 0 23644 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_251
timestamp 1644511149
transform 1 0 24196 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_98_253
timestamp 1644511149
transform 1 0 24380 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_98_265
timestamp 1644511149
transform 1 0 25484 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_98_269
timestamp 1644511149
transform 1 0 25852 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_98_291
timestamp 1644511149
transform 1 0 27876 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_98_303
timestamp 1644511149
transform 1 0 28980 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_98_307
timestamp 1644511149
transform 1 0 29348 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_98_309
timestamp 1644511149
transform 1 0 29532 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_321
timestamp 1644511149
transform 1 0 30636 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_333
timestamp 1644511149
transform 1 0 31740 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_98_345
timestamp 1644511149
transform 1 0 32844 0 1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_98_356
timestamp 1644511149
transform 1 0 33856 0 1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_98_365
timestamp 1644511149
transform 1 0 34684 0 1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_98_373
timestamp 1644511149
transform 1 0 35420 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_98_397
timestamp 1644511149
transform 1 0 37628 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_98_409
timestamp 1644511149
transform 1 0 38732 0 1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_98_417
timestamp 1644511149
transform 1 0 39468 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_98_421
timestamp 1644511149
transform 1 0 39836 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_98_433
timestamp 1644511149
transform 1 0 40940 0 1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_98_441
timestamp 1644511149
transform 1 0 41676 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_98_465
timestamp 1644511149
transform 1 0 43884 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_98_472
timestamp 1644511149
transform 1 0 44528 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_98_477
timestamp 1644511149
transform 1 0 44988 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_489
timestamp 1644511149
transform 1 0 46092 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_501
timestamp 1644511149
transform 1 0 47196 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_513
timestamp 1644511149
transform 1 0 48300 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_525
timestamp 1644511149
transform 1 0 49404 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_531
timestamp 1644511149
transform 1 0 49956 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_98_536
timestamp 1644511149
transform 1 0 50416 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_548
timestamp 1644511149
transform 1 0 51520 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_98_560
timestamp 1644511149
transform 1 0 52624 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_98_564
timestamp 1644511149
transform 1 0 52992 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_98_568
timestamp 1644511149
transform 1 0 53360 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_98_580
timestamp 1644511149
transform 1 0 54464 0 1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_98_589
timestamp 1644511149
transform 1 0 55292 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_601
timestamp 1644511149
transform 1 0 56396 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_613
timestamp 1644511149
transform 1 0 57500 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_3
timestamp 1644511149
transform 1 0 1380 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_15
timestamp 1644511149
transform 1 0 2484 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_27
timestamp 1644511149
transform 1 0 3588 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_39
timestamp 1644511149
transform 1 0 4692 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_99_51
timestamp 1644511149
transform 1 0 5796 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_99_55
timestamp 1644511149
transform 1 0 6164 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_99_57
timestamp 1644511149
transform 1 0 6348 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_99_81
timestamp 1644511149
transform 1 0 8556 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_99_106
timestamp 1644511149
transform 1 0 10856 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_99_113
timestamp 1644511149
transform 1 0 11500 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_125
timestamp 1644511149
transform 1 0 12604 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_137
timestamp 1644511149
transform 1 0 13708 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_149
timestamp 1644511149
transform 1 0 14812 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_161
timestamp 1644511149
transform 1 0 15916 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_167
timestamp 1644511149
transform 1 0 16468 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_99_169
timestamp 1644511149
transform 1 0 16652 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_181
timestamp 1644511149
transform 1 0 17756 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_193
timestamp 1644511149
transform 1 0 18860 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_205
timestamp 1644511149
transform 1 0 19964 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_217
timestamp 1644511149
transform 1 0 21068 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_223
timestamp 1644511149
transform 1 0 21620 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_99_225
timestamp 1644511149
transform 1 0 21804 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_237
timestamp 1644511149
transform 1 0 22908 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_249
timestamp 1644511149
transform 1 0 24012 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_261
timestamp 1644511149
transform 1 0 25116 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_273
timestamp 1644511149
transform 1 0 26220 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_279
timestamp 1644511149
transform 1 0 26772 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_99_281
timestamp 1644511149
transform 1 0 26956 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_293
timestamp 1644511149
transform 1 0 28060 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_305
timestamp 1644511149
transform 1 0 29164 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_317
timestamp 1644511149
transform 1 0 30268 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_329
timestamp 1644511149
transform 1 0 31372 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_335
timestamp 1644511149
transform 1 0 31924 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_99_337
timestamp 1644511149
transform 1 0 32108 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_99_349
timestamp 1644511149
transform 1 0 33212 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_99_373
timestamp 1644511149
transform 1 0 35420 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_385
timestamp 1644511149
transform 1 0 36524 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_391
timestamp 1644511149
transform 1 0 37076 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_99_393
timestamp 1644511149
transform 1 0 37260 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_405
timestamp 1644511149
transform 1 0 38364 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_417
timestamp 1644511149
transform 1 0 39468 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_429
timestamp 1644511149
transform 1 0 40572 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_441
timestamp 1644511149
transform 1 0 41676 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_447
timestamp 1644511149
transform 1 0 42228 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_99_452
timestamp 1644511149
transform 1 0 42688 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_99_479
timestamp 1644511149
transform 1 0 45172 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_491
timestamp 1644511149
transform 1 0 46276 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_99_503
timestamp 1644511149
transform 1 0 47380 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_99_505
timestamp 1644511149
transform 1 0 47564 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_517
timestamp 1644511149
transform 1 0 48668 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_99_529
timestamp 1644511149
transform 1 0 49772 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_99_551
timestamp 1644511149
transform 1 0 51796 0 -1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_99_559
timestamp 1644511149
transform 1 0 52532 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_99_561
timestamp 1644511149
transform 1 0 52716 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_99_583
timestamp 1644511149
transform 1 0 54740 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_595
timestamp 1644511149
transform 1 0 55844 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_99_607
timestamp 1644511149
transform 1 0 56948 0 -1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_99_615
timestamp 1644511149
transform 1 0 57684 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_99_617
timestamp 1644511149
transform 1 0 57868 0 -1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_100_3
timestamp 1644511149
transform 1 0 1380 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_15
timestamp 1644511149
transform 1 0 2484 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_100_27
timestamp 1644511149
transform 1 0 3588 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_100_29
timestamp 1644511149
transform 1 0 3772 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_41
timestamp 1644511149
transform 1 0 4876 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_53
timestamp 1644511149
transform 1 0 5980 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_65
timestamp 1644511149
transform 1 0 7084 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_100_74
timestamp 1644511149
transform 1 0 7912 0 1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_100_82
timestamp 1644511149
transform 1 0 8648 0 1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_100_85
timestamp 1644511149
transform 1 0 8924 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_100_89
timestamp 1644511149
transform 1 0 9292 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_101
timestamp 1644511149
transform 1 0 10396 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_113
timestamp 1644511149
transform 1 0 11500 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_125
timestamp 1644511149
transform 1 0 12604 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_100_137
timestamp 1644511149
transform 1 0 13708 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_100_141
timestamp 1644511149
transform 1 0 14076 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_153
timestamp 1644511149
transform 1 0 15180 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_165
timestamp 1644511149
transform 1 0 16284 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_177
timestamp 1644511149
transform 1 0 17388 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_189
timestamp 1644511149
transform 1 0 18492 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_195
timestamp 1644511149
transform 1 0 19044 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_100_197
timestamp 1644511149
transform 1 0 19228 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_209
timestamp 1644511149
transform 1 0 20332 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_221
timestamp 1644511149
transform 1 0 21436 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_233
timestamp 1644511149
transform 1 0 22540 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_245
timestamp 1644511149
transform 1 0 23644 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_251
timestamp 1644511149
transform 1 0 24196 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_100_253
timestamp 1644511149
transform 1 0 24380 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_265
timestamp 1644511149
transform 1 0 25484 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_100_274
timestamp 1644511149
transform 1 0 26312 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_286
timestamp 1644511149
transform 1 0 27416 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_100_298
timestamp 1644511149
transform 1 0 28520 0 1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_100_306
timestamp 1644511149
transform 1 0 29256 0 1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_100_309
timestamp 1644511149
transform 1 0 29532 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_321
timestamp 1644511149
transform 1 0 30636 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_333
timestamp 1644511149
transform 1 0 31740 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_100_345
timestamp 1644511149
transform 1 0 32844 0 1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_100_356
timestamp 1644511149
transform 1 0 33856 0 1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_100_365
timestamp 1644511149
transform 1 0 34684 0 1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_100_373
timestamp 1644511149
transform 1 0 35420 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_100_379
timestamp 1644511149
transform 1 0 35972 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_391
timestamp 1644511149
transform 1 0 37076 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_403
timestamp 1644511149
transform 1 0 38180 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_100_415
timestamp 1644511149
transform 1 0 39284 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_100_419
timestamp 1644511149
transform 1 0 39652 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_100_421
timestamp 1644511149
transform 1 0 39836 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_433
timestamp 1644511149
transform 1 0 40940 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_100_445
timestamp 1644511149
transform 1 0 42044 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_100_449
timestamp 1644511149
transform 1 0 42412 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_100_453
timestamp 1644511149
transform 1 0 42780 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_100_460
timestamp 1644511149
transform 1 0 43424 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_100_472
timestamp 1644511149
transform 1 0 44528 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_100_477
timestamp 1644511149
transform 1 0 44988 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_489
timestamp 1644511149
transform 1 0 46092 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_501
timestamp 1644511149
transform 1 0 47196 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_513
timestamp 1644511149
transform 1 0 48300 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_525
timestamp 1644511149
transform 1 0 49404 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_531
timestamp 1644511149
transform 1 0 49956 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_100_536
timestamp 1644511149
transform 1 0 50416 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_548
timestamp 1644511149
transform 1 0 51520 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_100_560
timestamp 1644511149
transform 1 0 52624 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_100_566
timestamp 1644511149
transform 1 0 53176 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_100_578
timestamp 1644511149
transform 1 0 54280 0 1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_100_586
timestamp 1644511149
transform 1 0 55016 0 1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_100_589
timestamp 1644511149
transform 1 0 55292 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_601
timestamp 1644511149
transform 1 0 56396 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_613
timestamp 1644511149
transform 1 0 57500 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_3
timestamp 1644511149
transform 1 0 1380 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_15
timestamp 1644511149
transform 1 0 2484 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_101_27
timestamp 1644511149
transform 1 0 3588 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_101_29
timestamp 1644511149
transform 1 0 3772 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_41
timestamp 1644511149
transform 1 0 4876 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_101_53
timestamp 1644511149
transform 1 0 5980 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_101_57
timestamp 1644511149
transform 1 0 6348 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_69
timestamp 1644511149
transform 1 0 7452 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_101_81
timestamp 1644511149
transform 1 0 8556 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_101_85
timestamp 1644511149
transform 1 0 8924 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_97
timestamp 1644511149
transform 1 0 10028 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_101_109
timestamp 1644511149
transform 1 0 11132 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_101_113
timestamp 1644511149
transform 1 0 11500 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_125
timestamp 1644511149
transform 1 0 12604 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_101_137
timestamp 1644511149
transform 1 0 13708 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_101_141
timestamp 1644511149
transform 1 0 14076 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_153
timestamp 1644511149
transform 1 0 15180 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_101_165
timestamp 1644511149
transform 1 0 16284 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_101_169
timestamp 1644511149
transform 1 0 16652 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_181
timestamp 1644511149
transform 1 0 17756 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_101_193
timestamp 1644511149
transform 1 0 18860 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_101_197
timestamp 1644511149
transform 1 0 19228 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_209
timestamp 1644511149
transform 1 0 20332 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_101_221
timestamp 1644511149
transform 1 0 21436 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_101_225
timestamp 1644511149
transform 1 0 21804 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_237
timestamp 1644511149
transform 1 0 22908 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_101_249
timestamp 1644511149
transform 1 0 24012 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_101_253
timestamp 1644511149
transform 1 0 24380 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_265
timestamp 1644511149
transform 1 0 25484 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_101_277
timestamp 1644511149
transform 1 0 26588 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_101_281
timestamp 1644511149
transform 1 0 26956 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_293
timestamp 1644511149
transform 1 0 28060 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_101_305
timestamp 1644511149
transform 1 0 29164 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_101_309
timestamp 1644511149
transform 1 0 29532 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_321
timestamp 1644511149
transform 1 0 30636 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_101_333
timestamp 1644511149
transform 1 0 31740 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_101_337
timestamp 1644511149
transform 1 0 32108 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_349
timestamp 1644511149
transform 1 0 33212 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_101_361
timestamp 1644511149
transform 1 0 34316 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_101_365
timestamp 1644511149
transform 1 0 34684 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_377
timestamp 1644511149
transform 1 0 35788 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_101_389
timestamp 1644511149
transform 1 0 36892 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_101_393
timestamp 1644511149
transform 1 0 37260 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_405
timestamp 1644511149
transform 1 0 38364 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_101_417
timestamp 1644511149
transform 1 0 39468 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_101_421
timestamp 1644511149
transform 1 0 39836 0 -1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_101_429
timestamp 1644511149
transform 1 0 40572 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_101_444
timestamp 1644511149
transform 1 0 41952 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_101_449
timestamp 1644511149
transform 1 0 42412 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_461
timestamp 1644511149
transform 1 0 43516 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_101_473
timestamp 1644511149
transform 1 0 44620 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_101_477
timestamp 1644511149
transform 1 0 44988 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_489
timestamp 1644511149
transform 1 0 46092 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_101_501
timestamp 1644511149
transform 1 0 47196 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_101_505
timestamp 1644511149
transform 1 0 47564 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_517
timestamp 1644511149
transform 1 0 48668 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_101_529
timestamp 1644511149
transform 1 0 49772 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_101_533
timestamp 1644511149
transform 1 0 50140 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_545
timestamp 1644511149
transform 1 0 51244 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_101_557
timestamp 1644511149
transform 1 0 52348 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_101_561
timestamp 1644511149
transform 1 0 52716 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_573
timestamp 1644511149
transform 1 0 53820 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_101_585
timestamp 1644511149
transform 1 0 54924 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_101_589
timestamp 1644511149
transform 1 0 55292 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_601
timestamp 1644511149
transform 1 0 56396 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_101_613
timestamp 1644511149
transform 1 0 57500 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_101_617
timestamp 1644511149
transform 1 0 57868 0 -1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1644511149
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1644511149
transform -1 0 58880 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1644511149
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1644511149
transform -1 0 58880 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1644511149
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1644511149
transform -1 0 58880 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1644511149
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1644511149
transform -1 0 58880 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1644511149
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1644511149
transform -1 0 58880 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1644511149
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1644511149
transform -1 0 58880 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1644511149
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1644511149
transform -1 0 58880 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1644511149
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1644511149
transform -1 0 58880 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1644511149
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1644511149
transform -1 0 58880 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1644511149
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1644511149
transform -1 0 58880 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1644511149
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1644511149
transform -1 0 58880 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1644511149
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1644511149
transform -1 0 58880 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1644511149
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1644511149
transform -1 0 58880 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1644511149
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1644511149
transform -1 0 58880 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1644511149
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1644511149
transform -1 0 58880 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1644511149
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1644511149
transform -1 0 58880 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1644511149
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1644511149
transform -1 0 58880 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1644511149
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1644511149
transform -1 0 58880 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1644511149
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1644511149
transform -1 0 58880 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1644511149
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1644511149
transform -1 0 58880 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1644511149
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1644511149
transform -1 0 58880 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1644511149
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1644511149
transform -1 0 58880 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1644511149
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1644511149
transform -1 0 58880 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1644511149
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1644511149
transform -1 0 58880 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1644511149
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1644511149
transform -1 0 58880 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1644511149
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1644511149
transform -1 0 58880 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1644511149
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1644511149
transform -1 0 58880 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1644511149
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1644511149
transform -1 0 58880 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1644511149
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1644511149
transform -1 0 58880 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1644511149
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1644511149
transform -1 0 58880 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1644511149
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1644511149
transform -1 0 58880 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1644511149
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1644511149
transform -1 0 58880 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1644511149
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1644511149
transform -1 0 58880 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1644511149
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1644511149
transform -1 0 58880 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1644511149
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1644511149
transform -1 0 58880 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1644511149
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1644511149
transform -1 0 58880 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1644511149
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1644511149
transform -1 0 58880 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1644511149
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1644511149
transform -1 0 58880 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1644511149
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1644511149
transform -1 0 58880 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1644511149
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1644511149
transform -1 0 58880 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1644511149
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1644511149
transform -1 0 58880 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1644511149
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1644511149
transform -1 0 58880 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1644511149
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1644511149
transform -1 0 58880 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1644511149
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1644511149
transform -1 0 58880 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1644511149
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1644511149
transform -1 0 58880 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1644511149
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1644511149
transform -1 0 58880 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1644511149
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1644511149
transform -1 0 58880 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1644511149
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1644511149
transform -1 0 58880 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1644511149
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1644511149
transform -1 0 58880 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1644511149
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1644511149
transform -1 0 58880 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1644511149
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1644511149
transform -1 0 58880 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1644511149
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1644511149
transform -1 0 58880 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1644511149
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1644511149
transform -1 0 58880 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1644511149
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1644511149
transform -1 0 58880 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1644511149
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1644511149
transform -1 0 58880 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1644511149
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1644511149
transform -1 0 58880 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1644511149
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1644511149
transform -1 0 58880 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1644511149
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1644511149
transform -1 0 58880 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 1644511149
transform 1 0 1104 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 1644511149
transform -1 0 58880 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 1644511149
transform 1 0 1104 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 1644511149
transform -1 0 58880 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 1644511149
transform 1 0 1104 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 1644511149
transform -1 0 58880 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_122
timestamp 1644511149
transform 1 0 1104 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_123
timestamp 1644511149
transform -1 0 58880 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_124
timestamp 1644511149
transform 1 0 1104 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_125
timestamp 1644511149
transform -1 0 58880 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_126
timestamp 1644511149
transform 1 0 1104 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_127
timestamp 1644511149
transform -1 0 58880 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_128
timestamp 1644511149
transform 1 0 1104 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_129
timestamp 1644511149
transform -1 0 58880 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_130
timestamp 1644511149
transform 1 0 1104 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_131
timestamp 1644511149
transform -1 0 58880 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_132
timestamp 1644511149
transform 1 0 1104 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_133
timestamp 1644511149
transform -1 0 58880 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_134
timestamp 1644511149
transform 1 0 1104 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_135
timestamp 1644511149
transform -1 0 58880 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_136
timestamp 1644511149
transform 1 0 1104 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_137
timestamp 1644511149
transform -1 0 58880 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_138
timestamp 1644511149
transform 1 0 1104 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_139
timestamp 1644511149
transform -1 0 58880 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_140
timestamp 1644511149
transform 1 0 1104 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_141
timestamp 1644511149
transform -1 0 58880 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_142
timestamp 1644511149
transform 1 0 1104 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_143
timestamp 1644511149
transform -1 0 58880 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_144
timestamp 1644511149
transform 1 0 1104 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_145
timestamp 1644511149
transform -1 0 58880 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_146
timestamp 1644511149
transform 1 0 1104 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_147
timestamp 1644511149
transform -1 0 58880 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_148
timestamp 1644511149
transform 1 0 1104 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_149
timestamp 1644511149
transform -1 0 58880 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_150
timestamp 1644511149
transform 1 0 1104 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_151
timestamp 1644511149
transform -1 0 58880 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_152
timestamp 1644511149
transform 1 0 1104 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_153
timestamp 1644511149
transform -1 0 58880 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_154
timestamp 1644511149
transform 1 0 1104 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_155
timestamp 1644511149
transform -1 0 58880 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_156
timestamp 1644511149
transform 1 0 1104 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_157
timestamp 1644511149
transform -1 0 58880 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_158
timestamp 1644511149
transform 1 0 1104 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_159
timestamp 1644511149
transform -1 0 58880 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_160
timestamp 1644511149
transform 1 0 1104 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_161
timestamp 1644511149
transform -1 0 58880 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_162
timestamp 1644511149
transform 1 0 1104 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_163
timestamp 1644511149
transform -1 0 58880 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_164
timestamp 1644511149
transform 1 0 1104 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_165
timestamp 1644511149
transform -1 0 58880 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_166
timestamp 1644511149
transform 1 0 1104 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_167
timestamp 1644511149
transform -1 0 58880 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_168
timestamp 1644511149
transform 1 0 1104 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_169
timestamp 1644511149
transform -1 0 58880 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_170
timestamp 1644511149
transform 1 0 1104 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_171
timestamp 1644511149
transform -1 0 58880 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_172
timestamp 1644511149
transform 1 0 1104 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_173
timestamp 1644511149
transform -1 0 58880 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_174
timestamp 1644511149
transform 1 0 1104 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_175
timestamp 1644511149
transform -1 0 58880 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_176
timestamp 1644511149
transform 1 0 1104 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_177
timestamp 1644511149
transform -1 0 58880 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_178
timestamp 1644511149
transform 1 0 1104 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_179
timestamp 1644511149
transform -1 0 58880 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_180
timestamp 1644511149
transform 1 0 1104 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_181
timestamp 1644511149
transform -1 0 58880 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_182
timestamp 1644511149
transform 1 0 1104 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_183
timestamp 1644511149
transform -1 0 58880 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_184
timestamp 1644511149
transform 1 0 1104 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_185
timestamp 1644511149
transform -1 0 58880 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_186
timestamp 1644511149
transform 1 0 1104 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_187
timestamp 1644511149
transform -1 0 58880 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_188
timestamp 1644511149
transform 1 0 1104 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_189
timestamp 1644511149
transform -1 0 58880 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_190
timestamp 1644511149
transform 1 0 1104 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_191
timestamp 1644511149
transform -1 0 58880 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_192
timestamp 1644511149
transform 1 0 1104 0 1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_193
timestamp 1644511149
transform -1 0 58880 0 1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_194
timestamp 1644511149
transform 1 0 1104 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_195
timestamp 1644511149
transform -1 0 58880 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_196
timestamp 1644511149
transform 1 0 1104 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_197
timestamp 1644511149
transform -1 0 58880 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_198
timestamp 1644511149
transform 1 0 1104 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_199
timestamp 1644511149
transform -1 0 58880 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_200
timestamp 1644511149
transform 1 0 1104 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_201
timestamp 1644511149
transform -1 0 58880 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_202
timestamp 1644511149
transform 1 0 1104 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_203
timestamp 1644511149
transform -1 0 58880 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1644511149
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1644511149
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1644511149
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1644511149
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1644511149
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1644511149
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1644511149
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1644511149
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1644511149
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1644511149
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1644511149
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1644511149
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1644511149
transform 1 0 37168 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1644511149
transform 1 0 39744 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1644511149
transform 1 0 42320 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1644511149
transform 1 0 44896 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1644511149
transform 1 0 47472 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1644511149
transform 1 0 50048 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1644511149
transform 1 0 52624 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1644511149
transform 1 0 55200 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1644511149
transform 1 0 57776 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1644511149
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1644511149
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1644511149
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1644511149
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1644511149
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1644511149
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1644511149
transform 1 0 37168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1644511149
transform 1 0 42320 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1644511149
transform 1 0 47472 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1644511149
transform 1 0 52624 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1644511149
transform 1 0 57776 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1644511149
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1644511149
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1644511149
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1644511149
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1644511149
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1644511149
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1644511149
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1644511149
transform 1 0 39744 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1644511149
transform 1 0 44896 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1644511149
transform 1 0 50048 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1644511149
transform 1 0 55200 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1644511149
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1644511149
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1644511149
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1644511149
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1644511149
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1644511149
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1644511149
transform 1 0 37168 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1644511149
transform 1 0 42320 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1644511149
transform 1 0 47472 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1644511149
transform 1 0 52624 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1644511149
transform 1 0 57776 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1644511149
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1644511149
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1644511149
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1644511149
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1644511149
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1644511149
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1644511149
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1644511149
transform 1 0 39744 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1644511149
transform 1 0 44896 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1644511149
transform 1 0 50048 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1644511149
transform 1 0 55200 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1644511149
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1644511149
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1644511149
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1644511149
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1644511149
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1644511149
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1644511149
transform 1 0 37168 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1644511149
transform 1 0 42320 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1644511149
transform 1 0 47472 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1644511149
transform 1 0 52624 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1644511149
transform 1 0 57776 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1644511149
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1644511149
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1644511149
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1644511149
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1644511149
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1644511149
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1644511149
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1644511149
transform 1 0 39744 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1644511149
transform 1 0 44896 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1644511149
transform 1 0 50048 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1644511149
transform 1 0 55200 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1644511149
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1644511149
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1644511149
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1644511149
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1644511149
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1644511149
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1644511149
transform 1 0 37168 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1644511149
transform 1 0 42320 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1644511149
transform 1 0 47472 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1644511149
transform 1 0 52624 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1644511149
transform 1 0 57776 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1644511149
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1644511149
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1644511149
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1644511149
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1644511149
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1644511149
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1644511149
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1644511149
transform 1 0 39744 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1644511149
transform 1 0 44896 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1644511149
transform 1 0 50048 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1644511149
transform 1 0 55200 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1644511149
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1644511149
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1644511149
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1644511149
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1644511149
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1644511149
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1644511149
transform 1 0 37168 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1644511149
transform 1 0 42320 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1644511149
transform 1 0 47472 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1644511149
transform 1 0 52624 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1644511149
transform 1 0 57776 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1644511149
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1644511149
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1644511149
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1644511149
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1644511149
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1644511149
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1644511149
transform 1 0 34592 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1644511149
transform 1 0 39744 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1644511149
transform 1 0 44896 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1644511149
transform 1 0 50048 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1644511149
transform 1 0 55200 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1644511149
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1644511149
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1644511149
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1644511149
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1644511149
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1644511149
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1644511149
transform 1 0 37168 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1644511149
transform 1 0 42320 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1644511149
transform 1 0 47472 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1644511149
transform 1 0 52624 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1644511149
transform 1 0 57776 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1644511149
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1644511149
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1644511149
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1644511149
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1644511149
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1644511149
transform 1 0 29440 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1644511149
transform 1 0 34592 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1644511149
transform 1 0 39744 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1644511149
transform 1 0 44896 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1644511149
transform 1 0 50048 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1644511149
transform 1 0 55200 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1644511149
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1644511149
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1644511149
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1644511149
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1644511149
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1644511149
transform 1 0 32016 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1644511149
transform 1 0 37168 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1644511149
transform 1 0 42320 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1644511149
transform 1 0 47472 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1644511149
transform 1 0 52624 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1644511149
transform 1 0 57776 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1644511149
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1644511149
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1644511149
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1644511149
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1644511149
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1644511149
transform 1 0 29440 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1644511149
transform 1 0 34592 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1644511149
transform 1 0 39744 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1644511149
transform 1 0 44896 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1644511149
transform 1 0 50048 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1644511149
transform 1 0 55200 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1644511149
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1644511149
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1644511149
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1644511149
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1644511149
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1644511149
transform 1 0 32016 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1644511149
transform 1 0 37168 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1644511149
transform 1 0 42320 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1644511149
transform 1 0 47472 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1644511149
transform 1 0 52624 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1644511149
transform 1 0 57776 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1644511149
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1644511149
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1644511149
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1644511149
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1644511149
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1644511149
transform 1 0 29440 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1644511149
transform 1 0 34592 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1644511149
transform 1 0 39744 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1644511149
transform 1 0 44896 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1644511149
transform 1 0 50048 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1644511149
transform 1 0 55200 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1644511149
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1644511149
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1644511149
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1644511149
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1644511149
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1644511149
transform 1 0 32016 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1644511149
transform 1 0 37168 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1644511149
transform 1 0 42320 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1644511149
transform 1 0 47472 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1644511149
transform 1 0 52624 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1644511149
transform 1 0 57776 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1644511149
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1644511149
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1644511149
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 1644511149
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 1644511149
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 1644511149
transform 1 0 29440 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 1644511149
transform 1 0 34592 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 1644511149
transform 1 0 39744 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_421
timestamp 1644511149
transform 1 0 44896 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_422
timestamp 1644511149
transform 1 0 50048 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_423
timestamp 1644511149
transform 1 0 55200 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_424
timestamp 1644511149
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_425
timestamp 1644511149
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_426
timestamp 1644511149
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_427
timestamp 1644511149
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_428
timestamp 1644511149
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_429
timestamp 1644511149
transform 1 0 32016 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_430
timestamp 1644511149
transform 1 0 37168 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_431
timestamp 1644511149
transform 1 0 42320 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_432
timestamp 1644511149
transform 1 0 47472 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_433
timestamp 1644511149
transform 1 0 52624 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_434
timestamp 1644511149
transform 1 0 57776 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_435
timestamp 1644511149
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_436
timestamp 1644511149
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_437
timestamp 1644511149
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_438
timestamp 1644511149
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_439
timestamp 1644511149
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_440
timestamp 1644511149
transform 1 0 29440 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_441
timestamp 1644511149
transform 1 0 34592 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_442
timestamp 1644511149
transform 1 0 39744 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_443
timestamp 1644511149
transform 1 0 44896 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_444
timestamp 1644511149
transform 1 0 50048 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_445
timestamp 1644511149
transform 1 0 55200 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_446
timestamp 1644511149
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_447
timestamp 1644511149
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_448
timestamp 1644511149
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_449
timestamp 1644511149
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_450
timestamp 1644511149
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_451
timestamp 1644511149
transform 1 0 32016 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_452
timestamp 1644511149
transform 1 0 37168 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_453
timestamp 1644511149
transform 1 0 42320 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_454
timestamp 1644511149
transform 1 0 47472 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_455
timestamp 1644511149
transform 1 0 52624 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_456
timestamp 1644511149
transform 1 0 57776 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_457
timestamp 1644511149
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_458
timestamp 1644511149
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_459
timestamp 1644511149
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_460
timestamp 1644511149
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_461
timestamp 1644511149
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_462
timestamp 1644511149
transform 1 0 29440 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_463
timestamp 1644511149
transform 1 0 34592 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_464
timestamp 1644511149
transform 1 0 39744 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_465
timestamp 1644511149
transform 1 0 44896 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_466
timestamp 1644511149
transform 1 0 50048 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_467
timestamp 1644511149
transform 1 0 55200 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_468
timestamp 1644511149
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_469
timestamp 1644511149
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_470
timestamp 1644511149
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_471
timestamp 1644511149
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_472
timestamp 1644511149
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_473
timestamp 1644511149
transform 1 0 32016 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_474
timestamp 1644511149
transform 1 0 37168 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_475
timestamp 1644511149
transform 1 0 42320 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_476
timestamp 1644511149
transform 1 0 47472 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_477
timestamp 1644511149
transform 1 0 52624 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_478
timestamp 1644511149
transform 1 0 57776 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_479
timestamp 1644511149
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_480
timestamp 1644511149
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_481
timestamp 1644511149
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_482
timestamp 1644511149
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_483
timestamp 1644511149
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_484
timestamp 1644511149
transform 1 0 29440 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_485
timestamp 1644511149
transform 1 0 34592 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_486
timestamp 1644511149
transform 1 0 39744 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_487
timestamp 1644511149
transform 1 0 44896 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_488
timestamp 1644511149
transform 1 0 50048 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_489
timestamp 1644511149
transform 1 0 55200 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_490
timestamp 1644511149
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_491
timestamp 1644511149
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_492
timestamp 1644511149
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_493
timestamp 1644511149
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_494
timestamp 1644511149
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_495
timestamp 1644511149
transform 1 0 32016 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_496
timestamp 1644511149
transform 1 0 37168 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_497
timestamp 1644511149
transform 1 0 42320 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_498
timestamp 1644511149
transform 1 0 47472 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_499
timestamp 1644511149
transform 1 0 52624 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_500
timestamp 1644511149
transform 1 0 57776 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_501
timestamp 1644511149
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_502
timestamp 1644511149
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_503
timestamp 1644511149
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_504
timestamp 1644511149
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_505
timestamp 1644511149
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_506
timestamp 1644511149
transform 1 0 29440 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_507
timestamp 1644511149
transform 1 0 34592 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_508
timestamp 1644511149
transform 1 0 39744 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_509
timestamp 1644511149
transform 1 0 44896 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_510
timestamp 1644511149
transform 1 0 50048 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_511
timestamp 1644511149
transform 1 0 55200 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_512
timestamp 1644511149
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_513
timestamp 1644511149
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_514
timestamp 1644511149
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_515
timestamp 1644511149
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_516
timestamp 1644511149
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_517
timestamp 1644511149
transform 1 0 32016 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_518
timestamp 1644511149
transform 1 0 37168 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_519
timestamp 1644511149
transform 1 0 42320 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_520
timestamp 1644511149
transform 1 0 47472 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_521
timestamp 1644511149
transform 1 0 52624 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_522
timestamp 1644511149
transform 1 0 57776 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_523
timestamp 1644511149
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_524
timestamp 1644511149
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_525
timestamp 1644511149
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_526
timestamp 1644511149
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_527
timestamp 1644511149
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_528
timestamp 1644511149
transform 1 0 29440 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_529
timestamp 1644511149
transform 1 0 34592 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_530
timestamp 1644511149
transform 1 0 39744 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_531
timestamp 1644511149
transform 1 0 44896 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_532
timestamp 1644511149
transform 1 0 50048 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_533
timestamp 1644511149
transform 1 0 55200 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_534
timestamp 1644511149
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_535
timestamp 1644511149
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_536
timestamp 1644511149
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_537
timestamp 1644511149
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_538
timestamp 1644511149
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_539
timestamp 1644511149
transform 1 0 32016 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_540
timestamp 1644511149
transform 1 0 37168 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_541
timestamp 1644511149
transform 1 0 42320 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_542
timestamp 1644511149
transform 1 0 47472 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_543
timestamp 1644511149
transform 1 0 52624 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_544
timestamp 1644511149
transform 1 0 57776 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_545
timestamp 1644511149
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_546
timestamp 1644511149
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_547
timestamp 1644511149
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_548
timestamp 1644511149
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_549
timestamp 1644511149
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_550
timestamp 1644511149
transform 1 0 29440 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_551
timestamp 1644511149
transform 1 0 34592 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_552
timestamp 1644511149
transform 1 0 39744 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_553
timestamp 1644511149
transform 1 0 44896 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_554
timestamp 1644511149
transform 1 0 50048 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_555
timestamp 1644511149
transform 1 0 55200 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_556
timestamp 1644511149
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_557
timestamp 1644511149
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_558
timestamp 1644511149
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_559
timestamp 1644511149
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_560
timestamp 1644511149
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_561
timestamp 1644511149
transform 1 0 32016 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_562
timestamp 1644511149
transform 1 0 37168 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_563
timestamp 1644511149
transform 1 0 42320 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_564
timestamp 1644511149
transform 1 0 47472 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_565
timestamp 1644511149
transform 1 0 52624 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_566
timestamp 1644511149
transform 1 0 57776 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_567
timestamp 1644511149
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_568
timestamp 1644511149
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_569
timestamp 1644511149
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_570
timestamp 1644511149
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_571
timestamp 1644511149
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_572
timestamp 1644511149
transform 1 0 29440 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_573
timestamp 1644511149
transform 1 0 34592 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_574
timestamp 1644511149
transform 1 0 39744 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_575
timestamp 1644511149
transform 1 0 44896 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_576
timestamp 1644511149
transform 1 0 50048 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_577
timestamp 1644511149
transform 1 0 55200 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_578
timestamp 1644511149
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_579
timestamp 1644511149
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_580
timestamp 1644511149
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_581
timestamp 1644511149
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_582
timestamp 1644511149
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_583
timestamp 1644511149
transform 1 0 32016 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_584
timestamp 1644511149
transform 1 0 37168 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_585
timestamp 1644511149
transform 1 0 42320 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_586
timestamp 1644511149
transform 1 0 47472 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_587
timestamp 1644511149
transform 1 0 52624 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_588
timestamp 1644511149
transform 1 0 57776 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_589
timestamp 1644511149
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_590
timestamp 1644511149
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_591
timestamp 1644511149
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_592
timestamp 1644511149
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_593
timestamp 1644511149
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_594
timestamp 1644511149
transform 1 0 29440 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_595
timestamp 1644511149
transform 1 0 34592 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_596
timestamp 1644511149
transform 1 0 39744 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_597
timestamp 1644511149
transform 1 0 44896 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_598
timestamp 1644511149
transform 1 0 50048 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_599
timestamp 1644511149
transform 1 0 55200 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_600
timestamp 1644511149
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_601
timestamp 1644511149
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_602
timestamp 1644511149
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_603
timestamp 1644511149
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_604
timestamp 1644511149
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_605
timestamp 1644511149
transform 1 0 32016 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_606
timestamp 1644511149
transform 1 0 37168 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_607
timestamp 1644511149
transform 1 0 42320 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_608
timestamp 1644511149
transform 1 0 47472 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_609
timestamp 1644511149
transform 1 0 52624 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_610
timestamp 1644511149
transform 1 0 57776 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_611
timestamp 1644511149
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_612
timestamp 1644511149
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_613
timestamp 1644511149
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_614
timestamp 1644511149
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_615
timestamp 1644511149
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_616
timestamp 1644511149
transform 1 0 29440 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_617
timestamp 1644511149
transform 1 0 34592 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_618
timestamp 1644511149
transform 1 0 39744 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_619
timestamp 1644511149
transform 1 0 44896 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_620
timestamp 1644511149
transform 1 0 50048 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_621
timestamp 1644511149
transform 1 0 55200 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_622
timestamp 1644511149
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_623
timestamp 1644511149
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_624
timestamp 1644511149
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_625
timestamp 1644511149
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_626
timestamp 1644511149
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_627
timestamp 1644511149
transform 1 0 32016 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_628
timestamp 1644511149
transform 1 0 37168 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_629
timestamp 1644511149
transform 1 0 42320 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_630
timestamp 1644511149
transform 1 0 47472 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_631
timestamp 1644511149
transform 1 0 52624 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_632
timestamp 1644511149
transform 1 0 57776 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_633
timestamp 1644511149
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_634
timestamp 1644511149
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_635
timestamp 1644511149
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_636
timestamp 1644511149
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_637
timestamp 1644511149
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_638
timestamp 1644511149
transform 1 0 29440 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_639
timestamp 1644511149
transform 1 0 34592 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_640
timestamp 1644511149
transform 1 0 39744 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_641
timestamp 1644511149
transform 1 0 44896 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_642
timestamp 1644511149
transform 1 0 50048 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_643
timestamp 1644511149
transform 1 0 55200 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_644
timestamp 1644511149
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_645
timestamp 1644511149
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_646
timestamp 1644511149
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_647
timestamp 1644511149
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_648
timestamp 1644511149
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_649
timestamp 1644511149
transform 1 0 32016 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_650
timestamp 1644511149
transform 1 0 37168 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_651
timestamp 1644511149
transform 1 0 42320 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_652
timestamp 1644511149
transform 1 0 47472 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_653
timestamp 1644511149
transform 1 0 52624 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_654
timestamp 1644511149
transform 1 0 57776 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_655
timestamp 1644511149
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_656
timestamp 1644511149
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_657
timestamp 1644511149
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_658
timestamp 1644511149
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_659
timestamp 1644511149
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_660
timestamp 1644511149
transform 1 0 29440 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_661
timestamp 1644511149
transform 1 0 34592 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_662
timestamp 1644511149
transform 1 0 39744 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_663
timestamp 1644511149
transform 1 0 44896 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_664
timestamp 1644511149
transform 1 0 50048 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_665
timestamp 1644511149
transform 1 0 55200 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_666
timestamp 1644511149
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_667
timestamp 1644511149
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_668
timestamp 1644511149
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_669
timestamp 1644511149
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_670
timestamp 1644511149
transform 1 0 26864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_671
timestamp 1644511149
transform 1 0 32016 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_672
timestamp 1644511149
transform 1 0 37168 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_673
timestamp 1644511149
transform 1 0 42320 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_674
timestamp 1644511149
transform 1 0 47472 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_675
timestamp 1644511149
transform 1 0 52624 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_676
timestamp 1644511149
transform 1 0 57776 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_677
timestamp 1644511149
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_678
timestamp 1644511149
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_679
timestamp 1644511149
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_680
timestamp 1644511149
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_681
timestamp 1644511149
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_682
timestamp 1644511149
transform 1 0 29440 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_683
timestamp 1644511149
transform 1 0 34592 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_684
timestamp 1644511149
transform 1 0 39744 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_685
timestamp 1644511149
transform 1 0 44896 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_686
timestamp 1644511149
transform 1 0 50048 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_687
timestamp 1644511149
transform 1 0 55200 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_688
timestamp 1644511149
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_689
timestamp 1644511149
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_690
timestamp 1644511149
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_691
timestamp 1644511149
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_692
timestamp 1644511149
transform 1 0 26864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_693
timestamp 1644511149
transform 1 0 32016 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_694
timestamp 1644511149
transform 1 0 37168 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_695
timestamp 1644511149
transform 1 0 42320 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_696
timestamp 1644511149
transform 1 0 47472 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_697
timestamp 1644511149
transform 1 0 52624 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_698
timestamp 1644511149
transform 1 0 57776 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_699
timestamp 1644511149
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_700
timestamp 1644511149
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_701
timestamp 1644511149
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_702
timestamp 1644511149
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_703
timestamp 1644511149
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_704
timestamp 1644511149
transform 1 0 29440 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_705
timestamp 1644511149
transform 1 0 34592 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_706
timestamp 1644511149
transform 1 0 39744 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_707
timestamp 1644511149
transform 1 0 44896 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_708
timestamp 1644511149
transform 1 0 50048 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_709
timestamp 1644511149
transform 1 0 55200 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_710
timestamp 1644511149
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_711
timestamp 1644511149
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_712
timestamp 1644511149
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_713
timestamp 1644511149
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_714
timestamp 1644511149
transform 1 0 26864 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_715
timestamp 1644511149
transform 1 0 32016 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_716
timestamp 1644511149
transform 1 0 37168 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_717
timestamp 1644511149
transform 1 0 42320 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_718
timestamp 1644511149
transform 1 0 47472 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_719
timestamp 1644511149
transform 1 0 52624 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_720
timestamp 1644511149
transform 1 0 57776 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_721
timestamp 1644511149
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_722
timestamp 1644511149
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_723
timestamp 1644511149
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_724
timestamp 1644511149
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_725
timestamp 1644511149
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_726
timestamp 1644511149
transform 1 0 29440 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_727
timestamp 1644511149
transform 1 0 34592 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_728
timestamp 1644511149
transform 1 0 39744 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_729
timestamp 1644511149
transform 1 0 44896 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_730
timestamp 1644511149
transform 1 0 50048 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_731
timestamp 1644511149
transform 1 0 55200 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_732
timestamp 1644511149
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_733
timestamp 1644511149
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_734
timestamp 1644511149
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_735
timestamp 1644511149
transform 1 0 21712 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_736
timestamp 1644511149
transform 1 0 26864 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_737
timestamp 1644511149
transform 1 0 32016 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_738
timestamp 1644511149
transform 1 0 37168 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_739
timestamp 1644511149
transform 1 0 42320 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_740
timestamp 1644511149
transform 1 0 47472 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_741
timestamp 1644511149
transform 1 0 52624 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_742
timestamp 1644511149
transform 1 0 57776 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_743
timestamp 1644511149
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_744
timestamp 1644511149
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_745
timestamp 1644511149
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_746
timestamp 1644511149
transform 1 0 19136 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_747
timestamp 1644511149
transform 1 0 24288 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_748
timestamp 1644511149
transform 1 0 29440 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_749
timestamp 1644511149
transform 1 0 34592 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_750
timestamp 1644511149
transform 1 0 39744 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_751
timestamp 1644511149
transform 1 0 44896 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_752
timestamp 1644511149
transform 1 0 50048 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_753
timestamp 1644511149
transform 1 0 55200 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_754
timestamp 1644511149
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_755
timestamp 1644511149
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_756
timestamp 1644511149
transform 1 0 16560 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_757
timestamp 1644511149
transform 1 0 21712 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_758
timestamp 1644511149
transform 1 0 26864 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_759
timestamp 1644511149
transform 1 0 32016 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_760
timestamp 1644511149
transform 1 0 37168 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_761
timestamp 1644511149
transform 1 0 42320 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_762
timestamp 1644511149
transform 1 0 47472 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_763
timestamp 1644511149
transform 1 0 52624 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_764
timestamp 1644511149
transform 1 0 57776 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_765
timestamp 1644511149
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_766
timestamp 1644511149
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_767
timestamp 1644511149
transform 1 0 13984 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_768
timestamp 1644511149
transform 1 0 19136 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_769
timestamp 1644511149
transform 1 0 24288 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_770
timestamp 1644511149
transform 1 0 29440 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_771
timestamp 1644511149
transform 1 0 34592 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_772
timestamp 1644511149
transform 1 0 39744 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_773
timestamp 1644511149
transform 1 0 44896 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_774
timestamp 1644511149
transform 1 0 50048 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_775
timestamp 1644511149
transform 1 0 55200 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_776
timestamp 1644511149
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_777
timestamp 1644511149
transform 1 0 11408 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_778
timestamp 1644511149
transform 1 0 16560 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_779
timestamp 1644511149
transform 1 0 21712 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_780
timestamp 1644511149
transform 1 0 26864 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_781
timestamp 1644511149
transform 1 0 32016 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_782
timestamp 1644511149
transform 1 0 37168 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_783
timestamp 1644511149
transform 1 0 42320 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_784
timestamp 1644511149
transform 1 0 47472 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_785
timestamp 1644511149
transform 1 0 52624 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_786
timestamp 1644511149
transform 1 0 57776 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_787
timestamp 1644511149
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_788
timestamp 1644511149
transform 1 0 8832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_789
timestamp 1644511149
transform 1 0 13984 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_790
timestamp 1644511149
transform 1 0 19136 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_791
timestamp 1644511149
transform 1 0 24288 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_792
timestamp 1644511149
transform 1 0 29440 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_793
timestamp 1644511149
transform 1 0 34592 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_794
timestamp 1644511149
transform 1 0 39744 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_795
timestamp 1644511149
transform 1 0 44896 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_796
timestamp 1644511149
transform 1 0 50048 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_797
timestamp 1644511149
transform 1 0 55200 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_798
timestamp 1644511149
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_799
timestamp 1644511149
transform 1 0 11408 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_800
timestamp 1644511149
transform 1 0 16560 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_801
timestamp 1644511149
transform 1 0 21712 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_802
timestamp 1644511149
transform 1 0 26864 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_803
timestamp 1644511149
transform 1 0 32016 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_804
timestamp 1644511149
transform 1 0 37168 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_805
timestamp 1644511149
transform 1 0 42320 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_806
timestamp 1644511149
transform 1 0 47472 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_807
timestamp 1644511149
transform 1 0 52624 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_808
timestamp 1644511149
transform 1 0 57776 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_809
timestamp 1644511149
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_810
timestamp 1644511149
transform 1 0 8832 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_811
timestamp 1644511149
transform 1 0 13984 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_812
timestamp 1644511149
transform 1 0 19136 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_813
timestamp 1644511149
transform 1 0 24288 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_814
timestamp 1644511149
transform 1 0 29440 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_815
timestamp 1644511149
transform 1 0 34592 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_816
timestamp 1644511149
transform 1 0 39744 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_817
timestamp 1644511149
transform 1 0 44896 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_818
timestamp 1644511149
transform 1 0 50048 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_819
timestamp 1644511149
transform 1 0 55200 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_820
timestamp 1644511149
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_821
timestamp 1644511149
transform 1 0 11408 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_822
timestamp 1644511149
transform 1 0 16560 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_823
timestamp 1644511149
transform 1 0 21712 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_824
timestamp 1644511149
transform 1 0 26864 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_825
timestamp 1644511149
transform 1 0 32016 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_826
timestamp 1644511149
transform 1 0 37168 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_827
timestamp 1644511149
transform 1 0 42320 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_828
timestamp 1644511149
transform 1 0 47472 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_829
timestamp 1644511149
transform 1 0 52624 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_830
timestamp 1644511149
transform 1 0 57776 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_831
timestamp 1644511149
transform 1 0 3680 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_832
timestamp 1644511149
transform 1 0 8832 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_833
timestamp 1644511149
transform 1 0 13984 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_834
timestamp 1644511149
transform 1 0 19136 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_835
timestamp 1644511149
transform 1 0 24288 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_836
timestamp 1644511149
transform 1 0 29440 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_837
timestamp 1644511149
transform 1 0 34592 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_838
timestamp 1644511149
transform 1 0 39744 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_839
timestamp 1644511149
transform 1 0 44896 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_840
timestamp 1644511149
transform 1 0 50048 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_841
timestamp 1644511149
transform 1 0 55200 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_842
timestamp 1644511149
transform 1 0 6256 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_843
timestamp 1644511149
transform 1 0 11408 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_844
timestamp 1644511149
transform 1 0 16560 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_845
timestamp 1644511149
transform 1 0 21712 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_846
timestamp 1644511149
transform 1 0 26864 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_847
timestamp 1644511149
transform 1 0 32016 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_848
timestamp 1644511149
transform 1 0 37168 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_849
timestamp 1644511149
transform 1 0 42320 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_850
timestamp 1644511149
transform 1 0 47472 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_851
timestamp 1644511149
transform 1 0 52624 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_852
timestamp 1644511149
transform 1 0 57776 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_853
timestamp 1644511149
transform 1 0 3680 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_854
timestamp 1644511149
transform 1 0 8832 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_855
timestamp 1644511149
transform 1 0 13984 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_856
timestamp 1644511149
transform 1 0 19136 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_857
timestamp 1644511149
transform 1 0 24288 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_858
timestamp 1644511149
transform 1 0 29440 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_859
timestamp 1644511149
transform 1 0 34592 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_860
timestamp 1644511149
transform 1 0 39744 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_861
timestamp 1644511149
transform 1 0 44896 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_862
timestamp 1644511149
transform 1 0 50048 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_863
timestamp 1644511149
transform 1 0 55200 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_864
timestamp 1644511149
transform 1 0 6256 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_865
timestamp 1644511149
transform 1 0 11408 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_866
timestamp 1644511149
transform 1 0 16560 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_867
timestamp 1644511149
transform 1 0 21712 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_868
timestamp 1644511149
transform 1 0 26864 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_869
timestamp 1644511149
transform 1 0 32016 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_870
timestamp 1644511149
transform 1 0 37168 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_871
timestamp 1644511149
transform 1 0 42320 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_872
timestamp 1644511149
transform 1 0 47472 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_873
timestamp 1644511149
transform 1 0 52624 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_874
timestamp 1644511149
transform 1 0 57776 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_875
timestamp 1644511149
transform 1 0 3680 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_876
timestamp 1644511149
transform 1 0 8832 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_877
timestamp 1644511149
transform 1 0 13984 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_878
timestamp 1644511149
transform 1 0 19136 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_879
timestamp 1644511149
transform 1 0 24288 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_880
timestamp 1644511149
transform 1 0 29440 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_881
timestamp 1644511149
transform 1 0 34592 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_882
timestamp 1644511149
transform 1 0 39744 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_883
timestamp 1644511149
transform 1 0 44896 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_884
timestamp 1644511149
transform 1 0 50048 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_885
timestamp 1644511149
transform 1 0 55200 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_886
timestamp 1644511149
transform 1 0 6256 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_887
timestamp 1644511149
transform 1 0 11408 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_888
timestamp 1644511149
transform 1 0 16560 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_889
timestamp 1644511149
transform 1 0 21712 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_890
timestamp 1644511149
transform 1 0 26864 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_891
timestamp 1644511149
transform 1 0 32016 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_892
timestamp 1644511149
transform 1 0 37168 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_893
timestamp 1644511149
transform 1 0 42320 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_894
timestamp 1644511149
transform 1 0 47472 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_895
timestamp 1644511149
transform 1 0 52624 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_896
timestamp 1644511149
transform 1 0 57776 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_897
timestamp 1644511149
transform 1 0 3680 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_898
timestamp 1644511149
transform 1 0 8832 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_899
timestamp 1644511149
transform 1 0 13984 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_900
timestamp 1644511149
transform 1 0 19136 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_901
timestamp 1644511149
transform 1 0 24288 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_902
timestamp 1644511149
transform 1 0 29440 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_903
timestamp 1644511149
transform 1 0 34592 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_904
timestamp 1644511149
transform 1 0 39744 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_905
timestamp 1644511149
transform 1 0 44896 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_906
timestamp 1644511149
transform 1 0 50048 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_907
timestamp 1644511149
transform 1 0 55200 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_908
timestamp 1644511149
transform 1 0 6256 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_909
timestamp 1644511149
transform 1 0 11408 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_910
timestamp 1644511149
transform 1 0 16560 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_911
timestamp 1644511149
transform 1 0 21712 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_912
timestamp 1644511149
transform 1 0 26864 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_913
timestamp 1644511149
transform 1 0 32016 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_914
timestamp 1644511149
transform 1 0 37168 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_915
timestamp 1644511149
transform 1 0 42320 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_916
timestamp 1644511149
transform 1 0 47472 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_917
timestamp 1644511149
transform 1 0 52624 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_918
timestamp 1644511149
transform 1 0 57776 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_919
timestamp 1644511149
transform 1 0 3680 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_920
timestamp 1644511149
transform 1 0 8832 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_921
timestamp 1644511149
transform 1 0 13984 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_922
timestamp 1644511149
transform 1 0 19136 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_923
timestamp 1644511149
transform 1 0 24288 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_924
timestamp 1644511149
transform 1 0 29440 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_925
timestamp 1644511149
transform 1 0 34592 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_926
timestamp 1644511149
transform 1 0 39744 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_927
timestamp 1644511149
transform 1 0 44896 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_928
timestamp 1644511149
transform 1 0 50048 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_929
timestamp 1644511149
transform 1 0 55200 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_930
timestamp 1644511149
transform 1 0 6256 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_931
timestamp 1644511149
transform 1 0 11408 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_932
timestamp 1644511149
transform 1 0 16560 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_933
timestamp 1644511149
transform 1 0 21712 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_934
timestamp 1644511149
transform 1 0 26864 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_935
timestamp 1644511149
transform 1 0 32016 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_936
timestamp 1644511149
transform 1 0 37168 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_937
timestamp 1644511149
transform 1 0 42320 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_938
timestamp 1644511149
transform 1 0 47472 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_939
timestamp 1644511149
transform 1 0 52624 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_940
timestamp 1644511149
transform 1 0 57776 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_941
timestamp 1644511149
transform 1 0 3680 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_942
timestamp 1644511149
transform 1 0 8832 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_943
timestamp 1644511149
transform 1 0 13984 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_944
timestamp 1644511149
transform 1 0 19136 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_945
timestamp 1644511149
transform 1 0 24288 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_946
timestamp 1644511149
transform 1 0 29440 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_947
timestamp 1644511149
transform 1 0 34592 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_948
timestamp 1644511149
transform 1 0 39744 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_949
timestamp 1644511149
transform 1 0 44896 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_950
timestamp 1644511149
transform 1 0 50048 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_951
timestamp 1644511149
transform 1 0 55200 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_952
timestamp 1644511149
transform 1 0 6256 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_953
timestamp 1644511149
transform 1 0 11408 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_954
timestamp 1644511149
transform 1 0 16560 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_955
timestamp 1644511149
transform 1 0 21712 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_956
timestamp 1644511149
transform 1 0 26864 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_957
timestamp 1644511149
transform 1 0 32016 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_958
timestamp 1644511149
transform 1 0 37168 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_959
timestamp 1644511149
transform 1 0 42320 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_960
timestamp 1644511149
transform 1 0 47472 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_961
timestamp 1644511149
transform 1 0 52624 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_962
timestamp 1644511149
transform 1 0 57776 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_963
timestamp 1644511149
transform 1 0 3680 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_964
timestamp 1644511149
transform 1 0 8832 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_965
timestamp 1644511149
transform 1 0 13984 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_966
timestamp 1644511149
transform 1 0 19136 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_967
timestamp 1644511149
transform 1 0 24288 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_968
timestamp 1644511149
transform 1 0 29440 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_969
timestamp 1644511149
transform 1 0 34592 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_970
timestamp 1644511149
transform 1 0 39744 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_971
timestamp 1644511149
transform 1 0 44896 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_972
timestamp 1644511149
transform 1 0 50048 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_973
timestamp 1644511149
transform 1 0 55200 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_974
timestamp 1644511149
transform 1 0 6256 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_975
timestamp 1644511149
transform 1 0 11408 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_976
timestamp 1644511149
transform 1 0 16560 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_977
timestamp 1644511149
transform 1 0 21712 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_978
timestamp 1644511149
transform 1 0 26864 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_979
timestamp 1644511149
transform 1 0 32016 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_980
timestamp 1644511149
transform 1 0 37168 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_981
timestamp 1644511149
transform 1 0 42320 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_982
timestamp 1644511149
transform 1 0 47472 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_983
timestamp 1644511149
transform 1 0 52624 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_984
timestamp 1644511149
transform 1 0 57776 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_985
timestamp 1644511149
transform 1 0 3680 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_986
timestamp 1644511149
transform 1 0 8832 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_987
timestamp 1644511149
transform 1 0 13984 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_988
timestamp 1644511149
transform 1 0 19136 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_989
timestamp 1644511149
transform 1 0 24288 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_990
timestamp 1644511149
transform 1 0 29440 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_991
timestamp 1644511149
transform 1 0 34592 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_992
timestamp 1644511149
transform 1 0 39744 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_993
timestamp 1644511149
transform 1 0 44896 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_994
timestamp 1644511149
transform 1 0 50048 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_995
timestamp 1644511149
transform 1 0 55200 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_996
timestamp 1644511149
transform 1 0 6256 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_997
timestamp 1644511149
transform 1 0 11408 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_998
timestamp 1644511149
transform 1 0 16560 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_999
timestamp 1644511149
transform 1 0 21712 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1000
timestamp 1644511149
transform 1 0 26864 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1001
timestamp 1644511149
transform 1 0 32016 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1002
timestamp 1644511149
transform 1 0 37168 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1003
timestamp 1644511149
transform 1 0 42320 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1004
timestamp 1644511149
transform 1 0 47472 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1005
timestamp 1644511149
transform 1 0 52624 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1006
timestamp 1644511149
transform 1 0 57776 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1007
timestamp 1644511149
transform 1 0 3680 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1008
timestamp 1644511149
transform 1 0 8832 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1009
timestamp 1644511149
transform 1 0 13984 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1010
timestamp 1644511149
transform 1 0 19136 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1011
timestamp 1644511149
transform 1 0 24288 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1012
timestamp 1644511149
transform 1 0 29440 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1013
timestamp 1644511149
transform 1 0 34592 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1014
timestamp 1644511149
transform 1 0 39744 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1015
timestamp 1644511149
transform 1 0 44896 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1016
timestamp 1644511149
transform 1 0 50048 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1017
timestamp 1644511149
transform 1 0 55200 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1018
timestamp 1644511149
transform 1 0 6256 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1019
timestamp 1644511149
transform 1 0 11408 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1020
timestamp 1644511149
transform 1 0 16560 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1021
timestamp 1644511149
transform 1 0 21712 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1022
timestamp 1644511149
transform 1 0 26864 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1023
timestamp 1644511149
transform 1 0 32016 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1024
timestamp 1644511149
transform 1 0 37168 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1025
timestamp 1644511149
transform 1 0 42320 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1026
timestamp 1644511149
transform 1 0 47472 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1027
timestamp 1644511149
transform 1 0 52624 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1028
timestamp 1644511149
transform 1 0 57776 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1029
timestamp 1644511149
transform 1 0 3680 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1030
timestamp 1644511149
transform 1 0 8832 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1031
timestamp 1644511149
transform 1 0 13984 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1032
timestamp 1644511149
transform 1 0 19136 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1033
timestamp 1644511149
transform 1 0 24288 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1034
timestamp 1644511149
transform 1 0 29440 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1035
timestamp 1644511149
transform 1 0 34592 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1036
timestamp 1644511149
transform 1 0 39744 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1037
timestamp 1644511149
transform 1 0 44896 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1038
timestamp 1644511149
transform 1 0 50048 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1039
timestamp 1644511149
transform 1 0 55200 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1040
timestamp 1644511149
transform 1 0 6256 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1041
timestamp 1644511149
transform 1 0 11408 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1042
timestamp 1644511149
transform 1 0 16560 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1043
timestamp 1644511149
transform 1 0 21712 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1044
timestamp 1644511149
transform 1 0 26864 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1045
timestamp 1644511149
transform 1 0 32016 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1046
timestamp 1644511149
transform 1 0 37168 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1047
timestamp 1644511149
transform 1 0 42320 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1048
timestamp 1644511149
transform 1 0 47472 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1049
timestamp 1644511149
transform 1 0 52624 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1050
timestamp 1644511149
transform 1 0 57776 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1051
timestamp 1644511149
transform 1 0 3680 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1052
timestamp 1644511149
transform 1 0 8832 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1053
timestamp 1644511149
transform 1 0 13984 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1054
timestamp 1644511149
transform 1 0 19136 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1055
timestamp 1644511149
transform 1 0 24288 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1056
timestamp 1644511149
transform 1 0 29440 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1057
timestamp 1644511149
transform 1 0 34592 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1058
timestamp 1644511149
transform 1 0 39744 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1059
timestamp 1644511149
transform 1 0 44896 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1060
timestamp 1644511149
transform 1 0 50048 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1061
timestamp 1644511149
transform 1 0 55200 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1062
timestamp 1644511149
transform 1 0 6256 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1063
timestamp 1644511149
transform 1 0 11408 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1064
timestamp 1644511149
transform 1 0 16560 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1065
timestamp 1644511149
transform 1 0 21712 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1066
timestamp 1644511149
transform 1 0 26864 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1067
timestamp 1644511149
transform 1 0 32016 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1068
timestamp 1644511149
transform 1 0 37168 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1069
timestamp 1644511149
transform 1 0 42320 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1070
timestamp 1644511149
transform 1 0 47472 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1071
timestamp 1644511149
transform 1 0 52624 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1072
timestamp 1644511149
transform 1 0 57776 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1073
timestamp 1644511149
transform 1 0 3680 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1074
timestamp 1644511149
transform 1 0 8832 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1075
timestamp 1644511149
transform 1 0 13984 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1076
timestamp 1644511149
transform 1 0 19136 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1077
timestamp 1644511149
transform 1 0 24288 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1078
timestamp 1644511149
transform 1 0 29440 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1079
timestamp 1644511149
transform 1 0 34592 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1080
timestamp 1644511149
transform 1 0 39744 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1081
timestamp 1644511149
transform 1 0 44896 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1082
timestamp 1644511149
transform 1 0 50048 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1083
timestamp 1644511149
transform 1 0 55200 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1084
timestamp 1644511149
transform 1 0 6256 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1085
timestamp 1644511149
transform 1 0 11408 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1086
timestamp 1644511149
transform 1 0 16560 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1087
timestamp 1644511149
transform 1 0 21712 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1088
timestamp 1644511149
transform 1 0 26864 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1089
timestamp 1644511149
transform 1 0 32016 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1090
timestamp 1644511149
transform 1 0 37168 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1091
timestamp 1644511149
transform 1 0 42320 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1092
timestamp 1644511149
transform 1 0 47472 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1093
timestamp 1644511149
transform 1 0 52624 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1094
timestamp 1644511149
transform 1 0 57776 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1095
timestamp 1644511149
transform 1 0 3680 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1096
timestamp 1644511149
transform 1 0 8832 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1097
timestamp 1644511149
transform 1 0 13984 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1098
timestamp 1644511149
transform 1 0 19136 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1099
timestamp 1644511149
transform 1 0 24288 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1100
timestamp 1644511149
transform 1 0 29440 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1101
timestamp 1644511149
transform 1 0 34592 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1102
timestamp 1644511149
transform 1 0 39744 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1103
timestamp 1644511149
transform 1 0 44896 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1104
timestamp 1644511149
transform 1 0 50048 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1105
timestamp 1644511149
transform 1 0 55200 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1106
timestamp 1644511149
transform 1 0 6256 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1107
timestamp 1644511149
transform 1 0 11408 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1108
timestamp 1644511149
transform 1 0 16560 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1109
timestamp 1644511149
transform 1 0 21712 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1110
timestamp 1644511149
transform 1 0 26864 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1111
timestamp 1644511149
transform 1 0 32016 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1112
timestamp 1644511149
transform 1 0 37168 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1113
timestamp 1644511149
transform 1 0 42320 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1114
timestamp 1644511149
transform 1 0 47472 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1115
timestamp 1644511149
transform 1 0 52624 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1116
timestamp 1644511149
transform 1 0 57776 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1117
timestamp 1644511149
transform 1 0 3680 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1118
timestamp 1644511149
transform 1 0 8832 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1119
timestamp 1644511149
transform 1 0 13984 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1120
timestamp 1644511149
transform 1 0 19136 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1121
timestamp 1644511149
transform 1 0 24288 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1122
timestamp 1644511149
transform 1 0 29440 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1123
timestamp 1644511149
transform 1 0 34592 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1124
timestamp 1644511149
transform 1 0 39744 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1125
timestamp 1644511149
transform 1 0 44896 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1126
timestamp 1644511149
transform 1 0 50048 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1127
timestamp 1644511149
transform 1 0 55200 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1128
timestamp 1644511149
transform 1 0 6256 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1129
timestamp 1644511149
transform 1 0 11408 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1130
timestamp 1644511149
transform 1 0 16560 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1131
timestamp 1644511149
transform 1 0 21712 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1132
timestamp 1644511149
transform 1 0 26864 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1133
timestamp 1644511149
transform 1 0 32016 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1134
timestamp 1644511149
transform 1 0 37168 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1135
timestamp 1644511149
transform 1 0 42320 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1136
timestamp 1644511149
transform 1 0 47472 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1137
timestamp 1644511149
transform 1 0 52624 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1138
timestamp 1644511149
transform 1 0 57776 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1139
timestamp 1644511149
transform 1 0 3680 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1140
timestamp 1644511149
transform 1 0 8832 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1141
timestamp 1644511149
transform 1 0 13984 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1142
timestamp 1644511149
transform 1 0 19136 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1143
timestamp 1644511149
transform 1 0 24288 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1144
timestamp 1644511149
transform 1 0 29440 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1145
timestamp 1644511149
transform 1 0 34592 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1146
timestamp 1644511149
transform 1 0 39744 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1147
timestamp 1644511149
transform 1 0 44896 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1148
timestamp 1644511149
transform 1 0 50048 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1149
timestamp 1644511149
transform 1 0 55200 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1150
timestamp 1644511149
transform 1 0 6256 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1151
timestamp 1644511149
transform 1 0 11408 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1152
timestamp 1644511149
transform 1 0 16560 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1153
timestamp 1644511149
transform 1 0 21712 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1154
timestamp 1644511149
transform 1 0 26864 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1155
timestamp 1644511149
transform 1 0 32016 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1156
timestamp 1644511149
transform 1 0 37168 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1157
timestamp 1644511149
transform 1 0 42320 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1158
timestamp 1644511149
transform 1 0 47472 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1159
timestamp 1644511149
transform 1 0 52624 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1160
timestamp 1644511149
transform 1 0 57776 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1161
timestamp 1644511149
transform 1 0 3680 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1162
timestamp 1644511149
transform 1 0 8832 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1163
timestamp 1644511149
transform 1 0 13984 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1164
timestamp 1644511149
transform 1 0 19136 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1165
timestamp 1644511149
transform 1 0 24288 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1166
timestamp 1644511149
transform 1 0 29440 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1167
timestamp 1644511149
transform 1 0 34592 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1168
timestamp 1644511149
transform 1 0 39744 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1169
timestamp 1644511149
transform 1 0 44896 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1170
timestamp 1644511149
transform 1 0 50048 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1171
timestamp 1644511149
transform 1 0 55200 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1172
timestamp 1644511149
transform 1 0 6256 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1173
timestamp 1644511149
transform 1 0 11408 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1174
timestamp 1644511149
transform 1 0 16560 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1175
timestamp 1644511149
transform 1 0 21712 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1176
timestamp 1644511149
transform 1 0 26864 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1177
timestamp 1644511149
transform 1 0 32016 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1178
timestamp 1644511149
transform 1 0 37168 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1179
timestamp 1644511149
transform 1 0 42320 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1180
timestamp 1644511149
transform 1 0 47472 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1181
timestamp 1644511149
transform 1 0 52624 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1182
timestamp 1644511149
transform 1 0 57776 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1183
timestamp 1644511149
transform 1 0 3680 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1184
timestamp 1644511149
transform 1 0 8832 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1185
timestamp 1644511149
transform 1 0 13984 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1186
timestamp 1644511149
transform 1 0 19136 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1187
timestamp 1644511149
transform 1 0 24288 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1188
timestamp 1644511149
transform 1 0 29440 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1189
timestamp 1644511149
transform 1 0 34592 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1190
timestamp 1644511149
transform 1 0 39744 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1191
timestamp 1644511149
transform 1 0 44896 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1192
timestamp 1644511149
transform 1 0 50048 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1193
timestamp 1644511149
transform 1 0 55200 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1194
timestamp 1644511149
transform 1 0 6256 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1195
timestamp 1644511149
transform 1 0 11408 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1196
timestamp 1644511149
transform 1 0 16560 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1197
timestamp 1644511149
transform 1 0 21712 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1198
timestamp 1644511149
transform 1 0 26864 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1199
timestamp 1644511149
transform 1 0 32016 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1200
timestamp 1644511149
transform 1 0 37168 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1201
timestamp 1644511149
transform 1 0 42320 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1202
timestamp 1644511149
transform 1 0 47472 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1203
timestamp 1644511149
transform 1 0 52624 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1204
timestamp 1644511149
transform 1 0 57776 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1205
timestamp 1644511149
transform 1 0 3680 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1206
timestamp 1644511149
transform 1 0 8832 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1207
timestamp 1644511149
transform 1 0 13984 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1208
timestamp 1644511149
transform 1 0 19136 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1209
timestamp 1644511149
transform 1 0 24288 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1210
timestamp 1644511149
transform 1 0 29440 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1211
timestamp 1644511149
transform 1 0 34592 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1212
timestamp 1644511149
transform 1 0 39744 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1213
timestamp 1644511149
transform 1 0 44896 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1214
timestamp 1644511149
transform 1 0 50048 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1215
timestamp 1644511149
transform 1 0 55200 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1216
timestamp 1644511149
transform 1 0 6256 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1217
timestamp 1644511149
transform 1 0 11408 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1218
timestamp 1644511149
transform 1 0 16560 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1219
timestamp 1644511149
transform 1 0 21712 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1220
timestamp 1644511149
transform 1 0 26864 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1221
timestamp 1644511149
transform 1 0 32016 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1222
timestamp 1644511149
transform 1 0 37168 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1223
timestamp 1644511149
transform 1 0 42320 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1224
timestamp 1644511149
transform 1 0 47472 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1225
timestamp 1644511149
transform 1 0 52624 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1226
timestamp 1644511149
transform 1 0 57776 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1227
timestamp 1644511149
transform 1 0 3680 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1228
timestamp 1644511149
transform 1 0 8832 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1229
timestamp 1644511149
transform 1 0 13984 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1230
timestamp 1644511149
transform 1 0 19136 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1231
timestamp 1644511149
transform 1 0 24288 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1232
timestamp 1644511149
transform 1 0 29440 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1233
timestamp 1644511149
transform 1 0 34592 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1234
timestamp 1644511149
transform 1 0 39744 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1235
timestamp 1644511149
transform 1 0 44896 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1236
timestamp 1644511149
transform 1 0 50048 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1237
timestamp 1644511149
transform 1 0 55200 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1238
timestamp 1644511149
transform 1 0 6256 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1239
timestamp 1644511149
transform 1 0 11408 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1240
timestamp 1644511149
transform 1 0 16560 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1241
timestamp 1644511149
transform 1 0 21712 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1242
timestamp 1644511149
transform 1 0 26864 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1243
timestamp 1644511149
transform 1 0 32016 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1244
timestamp 1644511149
transform 1 0 37168 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1245
timestamp 1644511149
transform 1 0 42320 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1246
timestamp 1644511149
transform 1 0 47472 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1247
timestamp 1644511149
transform 1 0 52624 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1248
timestamp 1644511149
transform 1 0 57776 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1249
timestamp 1644511149
transform 1 0 3680 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1250
timestamp 1644511149
transform 1 0 8832 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1251
timestamp 1644511149
transform 1 0 13984 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1252
timestamp 1644511149
transform 1 0 19136 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1253
timestamp 1644511149
transform 1 0 24288 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1254
timestamp 1644511149
transform 1 0 29440 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1255
timestamp 1644511149
transform 1 0 34592 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1256
timestamp 1644511149
transform 1 0 39744 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1257
timestamp 1644511149
transform 1 0 44896 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1258
timestamp 1644511149
transform 1 0 50048 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1259
timestamp 1644511149
transform 1 0 55200 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1260
timestamp 1644511149
transform 1 0 6256 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1261
timestamp 1644511149
transform 1 0 11408 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1262
timestamp 1644511149
transform 1 0 16560 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1263
timestamp 1644511149
transform 1 0 21712 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1264
timestamp 1644511149
transform 1 0 26864 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1265
timestamp 1644511149
transform 1 0 32016 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1266
timestamp 1644511149
transform 1 0 37168 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1267
timestamp 1644511149
transform 1 0 42320 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1268
timestamp 1644511149
transform 1 0 47472 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1269
timestamp 1644511149
transform 1 0 52624 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1270
timestamp 1644511149
transform 1 0 57776 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1271
timestamp 1644511149
transform 1 0 3680 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1272
timestamp 1644511149
transform 1 0 8832 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1273
timestamp 1644511149
transform 1 0 13984 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1274
timestamp 1644511149
transform 1 0 19136 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1275
timestamp 1644511149
transform 1 0 24288 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1276
timestamp 1644511149
transform 1 0 29440 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1277
timestamp 1644511149
transform 1 0 34592 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1278
timestamp 1644511149
transform 1 0 39744 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1279
timestamp 1644511149
transform 1 0 44896 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1280
timestamp 1644511149
transform 1 0 50048 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1281
timestamp 1644511149
transform 1 0 55200 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1282
timestamp 1644511149
transform 1 0 6256 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1283
timestamp 1644511149
transform 1 0 11408 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1284
timestamp 1644511149
transform 1 0 16560 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1285
timestamp 1644511149
transform 1 0 21712 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1286
timestamp 1644511149
transform 1 0 26864 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1287
timestamp 1644511149
transform 1 0 32016 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1288
timestamp 1644511149
transform 1 0 37168 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1289
timestamp 1644511149
transform 1 0 42320 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1290
timestamp 1644511149
transform 1 0 47472 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1291
timestamp 1644511149
transform 1 0 52624 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1292
timestamp 1644511149
transform 1 0 57776 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1293
timestamp 1644511149
transform 1 0 3680 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1294
timestamp 1644511149
transform 1 0 8832 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1295
timestamp 1644511149
transform 1 0 13984 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1296
timestamp 1644511149
transform 1 0 19136 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1297
timestamp 1644511149
transform 1 0 24288 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1298
timestamp 1644511149
transform 1 0 29440 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1299
timestamp 1644511149
transform 1 0 34592 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1300
timestamp 1644511149
transform 1 0 39744 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1301
timestamp 1644511149
transform 1 0 44896 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1302
timestamp 1644511149
transform 1 0 50048 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1303
timestamp 1644511149
transform 1 0 55200 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1304
timestamp 1644511149
transform 1 0 6256 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1305
timestamp 1644511149
transform 1 0 11408 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1306
timestamp 1644511149
transform 1 0 16560 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1307
timestamp 1644511149
transform 1 0 21712 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1308
timestamp 1644511149
transform 1 0 26864 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1309
timestamp 1644511149
transform 1 0 32016 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1310
timestamp 1644511149
transform 1 0 37168 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1311
timestamp 1644511149
transform 1 0 42320 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1312
timestamp 1644511149
transform 1 0 47472 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1313
timestamp 1644511149
transform 1 0 52624 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1314
timestamp 1644511149
transform 1 0 57776 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1315
timestamp 1644511149
transform 1 0 3680 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1316
timestamp 1644511149
transform 1 0 8832 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1317
timestamp 1644511149
transform 1 0 13984 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1318
timestamp 1644511149
transform 1 0 19136 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1319
timestamp 1644511149
transform 1 0 24288 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1320
timestamp 1644511149
transform 1 0 29440 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1321
timestamp 1644511149
transform 1 0 34592 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1322
timestamp 1644511149
transform 1 0 39744 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1323
timestamp 1644511149
transform 1 0 44896 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1324
timestamp 1644511149
transform 1 0 50048 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1325
timestamp 1644511149
transform 1 0 55200 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1326
timestamp 1644511149
transform 1 0 3680 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1327
timestamp 1644511149
transform 1 0 6256 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1328
timestamp 1644511149
transform 1 0 8832 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1329
timestamp 1644511149
transform 1 0 11408 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1330
timestamp 1644511149
transform 1 0 13984 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1331
timestamp 1644511149
transform 1 0 16560 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1332
timestamp 1644511149
transform 1 0 19136 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1333
timestamp 1644511149
transform 1 0 21712 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1334
timestamp 1644511149
transform 1 0 24288 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1335
timestamp 1644511149
transform 1 0 26864 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1336
timestamp 1644511149
transform 1 0 29440 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1337
timestamp 1644511149
transform 1 0 32016 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1338
timestamp 1644511149
transform 1 0 34592 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1339
timestamp 1644511149
transform 1 0 37168 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1340
timestamp 1644511149
transform 1 0 39744 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1341
timestamp 1644511149
transform 1 0 42320 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1342
timestamp 1644511149
transform 1 0 44896 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1343
timestamp 1644511149
transform 1 0 47472 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1344
timestamp 1644511149
transform 1 0 50048 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1345
timestamp 1644511149
transform 1 0 52624 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1346
timestamp 1644511149
transform 1 0 55200 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1347
timestamp 1644511149
transform 1 0 57776 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__buf_6  _237_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 7636 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_16  _238_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 57132 0 -1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__inv_2  _239_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 50416 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _240_
timestamp 1644511149
transform -1 0 15640 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _241_
timestamp 1644511149
transform 1 0 55660 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _242_
timestamp 1644511149
transform 1 0 54556 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _243_
timestamp 1644511149
transform 1 0 26036 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__buf_12  _244_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 8740 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_2  _245_
timestamp 1644511149
transform 1 0 33580 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _246_
timestamp 1644511149
transform -1 0 53360 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _247_
timestamp 1644511149
transform 1 0 57868 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _248_
timestamp 1644511149
transform -1 0 56948 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _249_
timestamp 1644511149
transform -1 0 4048 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__buf_8  _250_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 55384 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _251_
timestamp 1644511149
transform -1 0 44528 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _252_
timestamp 1644511149
transform 1 0 20700 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _253_
timestamp 1644511149
transform 1 0 35788 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _254_
timestamp 1644511149
transform 1 0 56304 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _255_
timestamp 1644511149
transform -1 0 18584 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_16  _256_
timestamp 1644511149
transform 1 0 7544 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__inv_2  _257_
timestamp 1644511149
transform 1 0 56948 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _258_
timestamp 1644511149
transform 1 0 56948 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _259_
timestamp 1644511149
transform -1 0 2576 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _260_
timestamp 1644511149
transform -1 0 2576 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _261_
timestamp 1644511149
transform -1 0 2576 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__buf_8  _262_
timestamp 1644511149
transform 1 0 7360 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _263_
timestamp 1644511149
transform -1 0 2576 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _264_
timestamp 1644511149
transform -1 0 2576 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _265_
timestamp 1644511149
transform 1 0 56764 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _266_
timestamp 1644511149
transform 1 0 44252 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _267_
timestamp 1644511149
transform -1 0 2576 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__buf_12  _268_
timestamp 1644511149
transform 1 0 7544 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_2  _269_
timestamp 1644511149
transform 1 0 9016 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _270_
timestamp 1644511149
transform 1 0 56304 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _271_
timestamp 1644511149
transform 1 0 51520 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _272_
timestamp 1644511149
transform -1 0 4048 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _273_
timestamp 1644511149
transform 1 0 4140 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _274_
timestamp 1644511149
transform -1 0 8372 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _275_
timestamp 1644511149
transform -1 0 57132 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _276_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 52716 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__nor3_1  _277_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 53084 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__and3b_1  _278_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 53360 0 -1 45696
box -38 -48 682 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _279_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 52716 0 1 45696
box -38 -48 958 592
use sky130_fd_sc_hd__and3b_1  _280_
timestamp 1644511149
transform -1 0 53360 0 -1 46784
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _281_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 50968 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _282_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 46460 0 1 51136
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _283_
timestamp 1644511149
transform -1 0 47840 0 1 51136
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _284_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 44712 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _285_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 46092 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _286_
timestamp 1644511149
transform -1 0 45264 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _287_
timestamp 1644511149
transform 1 0 46828 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _288_
timestamp 1644511149
transform -1 0 47012 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _289_
timestamp 1644511149
transform -1 0 46092 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _290_
timestamp 1644511149
transform -1 0 48668 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _291_
timestamp 1644511149
transform -1 0 49312 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _292_
timestamp 1644511149
transform -1 0 46828 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__and4bb_1  _293_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 50140 0 -1 52224
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _294_
timestamp 1644511149
transform 1 0 49220 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_1  _295_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 51152 0 -1 52224
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _296_
timestamp 1644511149
transform -1 0 50508 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__and4bb_1  _297_
timestamp 1644511149
transform 1 0 50140 0 1 52224
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _298_
timestamp 1644511149
transform -1 0 50876 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__and4bb_1  _299_
timestamp 1644511149
transform 1 0 49680 0 -1 53312
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _300_
timestamp 1644511149
transform -1 0 51796 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _301_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 47564 0 -1 52224
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_1  _302_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 47656 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _303_
timestamp 1644511149
transform 1 0 48208 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _304_
timestamp 1644511149
transform -1 0 45632 0 -1 43520
box -38 -48 958 592
use sky130_fd_sc_hd__inv_2  _305_
timestamp 1644511149
transform -1 0 46828 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _306_
timestamp 1644511149
transform 1 0 44620 0 -1 44608
box -38 -48 958 592
use sky130_fd_sc_hd__o211a_1  _307_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 47012 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _308_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 46552 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__or4b_1  _309_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 48116 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__o31ai_1  _310_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 46460 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _311_
timestamp 1644511149
transform 1 0 38088 0 1 45696
box -38 -48 958 592
use sky130_fd_sc_hd__nor2_1  _312_
timestamp 1644511149
transform 1 0 36524 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _313_
timestamp 1644511149
transform 1 0 37996 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _314_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 37076 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _315_
timestamp 1644511149
transform -1 0 37812 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _316_
timestamp 1644511149
transform 1 0 39284 0 -1 44608
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _317_
timestamp 1644511149
transform 1 0 39836 0 1 46784
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _318_
timestamp 1644511149
transform 1 0 37444 0 -1 47872
box -38 -48 958 592
use sky130_fd_sc_hd__nor3_1  _319_
timestamp 1644511149
transform -1 0 37076 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _320_
timestamp 1644511149
transform -1 0 37628 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _321_
timestamp 1644511149
transform 1 0 37260 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _322_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 38916 0 1 46784
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _323_
timestamp 1644511149
transform 1 0 39836 0 1 47872
box -38 -48 958 592
use sky130_fd_sc_hd__a21oi_1  _324_
timestamp 1644511149
transform 1 0 38180 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__a211oi_1  _325_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 36800 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _326_
timestamp 1644511149
transform -1 0 37536 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _327_
timestamp 1644511149
transform -1 0 37996 0 -1 48960
box -38 -48 498 592
use sky130_fd_sc_hd__nor3_1  _328_
timestamp 1644511149
transform -1 0 36800 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _329_
timestamp 1644511149
transform -1 0 39744 0 -1 50048
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _330_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 38364 0 -1 48960
box -38 -48 682 592
use sky130_fd_sc_hd__o21ba_1  _331_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 37904 0 -1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__a41o_1  _332_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 39376 0 -1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _333_
timestamp 1644511149
transform 1 0 39836 0 1 48960
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _334_
timestamp 1644511149
transform 1 0 38824 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _335_
timestamp 1644511149
transform -1 0 40756 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _336_
timestamp 1644511149
transform -1 0 44436 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _337_
timestamp 1644511149
transform 1 0 43700 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _338_
timestamp 1644511149
transform 1 0 43884 0 -1 43520
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _339_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 44068 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__or4_2  _340_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 46644 0 -1 43520
box -38 -48 682 592
use sky130_fd_sc_hd__o21bai_2  _341_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 45080 0 -1 45696
box -38 -48 866 592
use sky130_fd_sc_hd__a21oi_1  _342_
timestamp 1644511149
transform 1 0 43976 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _343_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 45448 0 1 42432
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _344_
timestamp 1644511149
transform 1 0 44988 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _345_
timestamp 1644511149
transform 1 0 44804 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _346_
timestamp 1644511149
transform 1 0 45540 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _347_
timestamp 1644511149
transform -1 0 46184 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _348_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 45908 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _349_
timestamp 1644511149
transform 1 0 46276 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _350_
timestamp 1644511149
transform 1 0 45448 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _351_
timestamp 1644511149
transform 1 0 49312 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__nor3_1  _352_
timestamp 1644511149
transform -1 0 48116 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__and2b_1  _353_
timestamp 1644511149
transform -1 0 49128 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _354_
timestamp 1644511149
transform 1 0 47472 0 1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _355_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 37260 0 -1 43520
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _356_
timestamp 1644511149
transform 1 0 36616 0 1 42432
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _357_
timestamp 1644511149
transform 1 0 37260 0 -1 44608
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _358_
timestamp 1644511149
transform 1 0 36248 0 1 45696
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _359_
timestamp 1644511149
transform 1 0 36340 0 1 46784
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _360_
timestamp 1644511149
transform 1 0 36248 0 1 48960
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _361_
timestamp 1644511149
transform 1 0 37536 0 1 50048
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _362_
timestamp 1644511149
transform 1 0 40480 0 -1 50048
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _363_
timestamp 1644511149
transform 1 0 43056 0 1 44608
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _364_
timestamp 1644511149
transform 1 0 43056 0 1 42432
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _365_
timestamp 1644511149
transform 1 0 45540 0 -1 42432
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _366_
timestamp 1644511149
transform 1 0 45724 0 1 41344
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _367_
timestamp 1644511149
transform 1 0 45632 0 1 45696
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _368_
timestamp 1644511149
transform -1 0 46920 0 -1 53312
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _369_
timestamp 1644511149
transform 1 0 44988 0 1 52224
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _370_
timestamp 1644511149
transform 1 0 47472 0 1 52224
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _371_
timestamp 1644511149
transform 1 0 47564 0 -1 50048
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _418__6 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 35972 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _419__7
timestamp 1644511149
transform 1 0 17204 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _420__8
timestamp 1644511149
transform -1 0 57500 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _421__9
timestamp 1644511149
transform -1 0 2300 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _422__10
timestamp 1644511149
transform -1 0 2300 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _423__11
timestamp 1644511149
transform -1 0 58144 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _424__12
timestamp 1644511149
transform -1 0 9292 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _425__13
timestamp 1644511149
transform -1 0 58144 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _426__14
timestamp 1644511149
transform 1 0 2208 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _427__15
timestamp 1644511149
transform -1 0 50416 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _428__16
timestamp 1644511149
transform -1 0 14720 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _429__17
timestamp 1644511149
transform -1 0 58144 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _430__18
timestamp 1644511149
transform -1 0 54740 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _431__19
timestamp 1644511149
transform -1 0 26312 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _432__20
timestamp 1644511149
transform -1 0 33856 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _433__21
timestamp 1644511149
transform -1 0 53176 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _434__22
timestamp 1644511149
transform 1 0 56580 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _435__23
timestamp 1644511149
transform -1 0 57500 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _436__24
timestamp 1644511149
transform 1 0 2392 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _437__25
timestamp 1644511149
transform -1 0 20976 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _438__26
timestamp 1644511149
transform -1 0 58144 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _439__27
timestamp 1644511149
transform 1 0 57868 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _440__28
timestamp 1644511149
transform -1 0 2300 0 1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _441__29
timestamp 1644511149
transform -1 0 2300 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _442__30
timestamp 1644511149
transform -1 0 2300 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _443__31
timestamp 1644511149
transform 1 0 44436 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _444__32
timestamp 1644511149
transform -1 0 2300 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _445__33
timestamp 1644511149
transform 1 0 7636 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _446__34
timestamp 1644511149
transform -1 0 4508 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _447__35
timestamp 1644511149
transform -1 0 51796 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _448__36
timestamp 1644511149
transform -1 0 58144 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _488__37
timestamp 1644511149
transform 1 0 42780 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _490__38
timestamp 1644511149
transform 1 0 41216 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _492__39
timestamp 1644511149
transform -1 0 44436 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _494__40
timestamp 1644511149
transform 1 0 42412 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _496__41
timestamp 1644511149
transform 1 0 42412 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _498__42
timestamp 1644511149
transform -1 0 42780 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _500__43
timestamp 1644511149
transform -1 0 43424 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _502_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 45172 0 -1 56576
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _503_
timestamp 1644511149
transform 1 0 35696 0 1 55488
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _504_
timestamp 1644511149
transform -1 0 18768 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _505_
timestamp 1644511149
transform 1 0 56304 0 1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _506_
timestamp 1644511149
transform 1 0 1932 0 -1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _507_
timestamp 1644511149
transform 1 0 1932 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _508_
timestamp 1644511149
transform 1 0 56304 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _509_
timestamp 1644511149
transform 1 0 8924 0 -1 56576
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _510_
timestamp 1644511149
transform 1 0 56304 0 1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _511_
timestamp 1644511149
transform -1 0 4048 0 -1 34816
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _512_
timestamp 1644511149
transform 1 0 49864 0 -1 56576
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _513_
timestamp 1644511149
transform 1 0 14444 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _514_
timestamp 1644511149
transform 1 0 56304 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _515_
timestamp 1644511149
transform 1 0 54464 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _516_
timestamp 1644511149
transform 1 0 25944 0 1 55488
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _517_
timestamp 1644511149
transform 1 0 33488 0 -1 56576
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _518_
timestamp 1644511149
transform 1 0 52808 0 -1 56576
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _519_
timestamp 1644511149
transform -1 0 57408 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _520_
timestamp 1644511149
transform 1 0 56304 0 1 41344
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _521_
timestamp 1644511149
transform -1 0 4232 0 -1 42432
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _522_
timestamp 1644511149
transform 1 0 20608 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _523_
timestamp 1644511149
transform 1 0 56304 0 1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _524_
timestamp 1644511149
transform -1 0 58236 0 1 28288
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _525_
timestamp 1644511149
transform 1 0 1932 0 -1 54400
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _526_
timestamp 1644511149
transform 1 0 1932 0 -1 47872
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _527_
timestamp 1644511149
transform 1 0 1932 0 -1 44608
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _528_
timestamp 1644511149
transform 1 0 44988 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _529_
timestamp 1644511149
transform 1 0 1932 0 -1 50048
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _530_
timestamp 1644511149
transform -1 0 8556 0 -1 56576
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _531_
timestamp 1644511149
transform 1 0 4048 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _532_
timestamp 1644511149
transform 1 0 51520 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _533_
timestamp 1644511149
transform 1 0 56304 0 1 23936
box -38 -48 1970 592
use sky130_fd_sc_hd__clkbuf_4  input1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 7176 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_8  input2
timestamp 1644511149
transform 1 0 40848 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1644511149
transform 1 0 57960 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__buf_12  input4
timestamp 1644511149
transform -1 0 58236 0 1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_6  input5
timestamp 1644511149
transform 1 0 24380 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__dlxtp_1  scan_wrapper_lesson1.latch\[0\] $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 50784 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  scan_wrapper_lesson1.latch\[1\]
timestamp 1644511149
transform 1 0 51060 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  scan_wrapper_lesson1.latch\[2\]
timestamp 1644511149
transform 1 0 50416 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  scan_wrapper_lesson1.latch\[3\]
timestamp 1644511149
transform 1 0 51888 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  scan_wrapper_lesson1.latch\[4\]
timestamp 1644511149
transform 1 0 51704 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  scan_wrapper_lesson1.latch\[5\]
timestamp 1644511149
transform 1 0 51060 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  scan_wrapper_lesson1.latch\[6\]
timestamp 1644511149
transform 1 0 50324 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  scan_wrapper_lesson1.latch\[7\]
timestamp 1644511149
transform 1 0 52716 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__sdfxtp_1  scan_wrapper_lesson1.scan_flop\[0\] $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 52256 0 1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__sdfxtp_1  scan_wrapper_lesson1.scan_flop\[1\]
timestamp 1644511149
transform -1 0 50876 0 -1 45696
box -38 -48 1970 592
use sky130_fd_sc_hd__sdfxtp_1  scan_wrapper_lesson1.scan_flop\[2\]
timestamp 1644511149
transform 1 0 47748 0 1 45696
box -38 -48 1970 592
use sky130_fd_sc_hd__sdfxtp_1  scan_wrapper_lesson1.scan_flop\[3\]
timestamp 1644511149
transform 1 0 49128 0 -1 44608
box -38 -48 1970 592
use sky130_fd_sc_hd__sdfxtp_1  scan_wrapper_lesson1.scan_flop\[4\]
timestamp 1644511149
transform 1 0 51796 0 1 42432
box -38 -48 1970 592
use sky130_fd_sc_hd__sdfxtp_1  scan_wrapper_lesson1.scan_flop\[5\]
timestamp 1644511149
transform -1 0 50324 0 -1 42432
box -38 -48 1970 592
use sky130_fd_sc_hd__sdfxtp_1  scan_wrapper_lesson1.scan_flop\[6\]
timestamp 1644511149
transform 1 0 47748 0 1 42432
box -38 -48 1970 592
use sky130_fd_sc_hd__sdfxtp_1  scan_wrapper_lesson1.scan_flop\[7\]
timestamp 1644511149
transform -1 0 50140 0 -1 43520
box -38 -48 1970 592
use sky130_fd_sc_hd__dlxtp_1  scan_wrapper_lesson2.latch\[0\]
timestamp 1644511149
transform -1 0 41584 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  scan_wrapper_lesson2.latch\[1\]
timestamp 1644511149
transform -1 0 41216 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__sdfxtp_1  scan_wrapper_lesson2.scan_flop\[0\]
timestamp 1644511149
transform -1 0 41952 0 1 42432
box -38 -48 1970 592
use sky130_fd_sc_hd__sdfxtp_1  scan_wrapper_lesson2.scan_flop\[1\]
timestamp 1644511149
transform 1 0 39836 0 -1 43520
box -38 -48 1970 592
use sky130_fd_sc_hd__sdfxtp_1  scan_wrapper_lesson2.scan_flop\[2\]
timestamp 1644511149
transform 1 0 39836 0 1 44608
box -38 -48 1970 592
use sky130_fd_sc_hd__sdfxtp_1  scan_wrapper_lesson2.scan_flop\[3\]
timestamp 1644511149
transform 1 0 39928 0 -1 45696
box -38 -48 1970 592
use sky130_fd_sc_hd__sdfxtp_1  scan_wrapper_lesson2.scan_flop\[4\]
timestamp 1644511149
transform 1 0 40020 0 -1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__sdfxtp_1  scan_wrapper_lesson2.scan_flop\[5\]
timestamp 1644511149
transform 1 0 40020 0 -1 47872
box -38 -48 1970 592
use sky130_fd_sc_hd__sdfxtp_1  scan_wrapper_lesson2.scan_flop\[6\]
timestamp 1644511149
transform 1 0 40848 0 1 48960
box -38 -48 1970 592
use sky130_fd_sc_hd__sdfxtp_1  scan_wrapper_lesson2.scan_flop\[7\]
timestamp 1644511149
transform 1 0 42412 0 -1 48960
box -38 -48 1970 592
use sky130_fd_sc_hd__dlxtp_1  scan_wrapper_lesson3.latch\[0\]
timestamp 1644511149
transform 1 0 44712 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  scan_wrapper_lesson3.latch\[1\]
timestamp 1644511149
transform -1 0 46736 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__sdfxtp_1  scan_wrapper_lesson3.scan_flop\[0\]
timestamp 1644511149
transform 1 0 43240 0 -1 50048
box -38 -48 1970 592
use sky130_fd_sc_hd__sdfxtp_1  scan_wrapper_lesson3.scan_flop\[1\]
timestamp 1644511149
transform 1 0 44988 0 1 48960
box -38 -48 1970 592
use sky130_fd_sc_hd__sdfxtp_1  scan_wrapper_lesson3.scan_flop\[2\]
timestamp 1644511149
transform 1 0 45724 0 1 47872
box -38 -48 1970 592
use sky130_fd_sc_hd__sdfxtp_1  scan_wrapper_lesson3.scan_flop\[3\]
timestamp 1644511149
transform 1 0 48576 0 -1 48960
box -38 -48 1970 592
use sky130_fd_sc_hd__sdfxtp_1  scan_wrapper_lesson3.scan_flop\[4\]
timestamp 1644511149
transform 1 0 50140 0 1 48960
box -38 -48 1970 592
use sky130_fd_sc_hd__sdfxtp_1  scan_wrapper_lesson3.scan_flop\[5\]
timestamp 1644511149
transform 1 0 50324 0 -1 50048
box -38 -48 1970 592
use sky130_fd_sc_hd__sdfxtp_1  scan_wrapper_lesson3.scan_flop\[6\]
timestamp 1644511149
transform 1 0 52440 0 1 48960
box -38 -48 1970 592
use sky130_fd_sc_hd__sdfxtp_1  scan_wrapper_lesson3.scan_flop\[7\]
timestamp 1644511149
transform 1 0 47748 0 1 48960
box -38 -48 1970 592
use sky130_fd_sc_hd__dlxtp_1  scan_wrapper_lesson4.latch\[0\]
timestamp 1644511149
transform -1 0 44528 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  scan_wrapper_lesson4.latch\[1\]
timestamp 1644511149
transform 1 0 43424 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__sdfxtp_1  scan_wrapper_lesson4.scan_flop\[0\]
timestamp 1644511149
transform -1 0 49496 0 -1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__sdfxtp_1  scan_wrapper_lesson4.scan_flop\[1\]
timestamp 1644511149
transform 1 0 42596 0 -1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__sdfxtp_1  scan_wrapper_lesson4.scan_flop\[2\]
timestamp 1644511149
transform -1 0 44344 0 -1 52224
box -38 -48 1970 592
use sky130_fd_sc_hd__sdfxtp_1  scan_wrapper_lesson4.scan_flop\[3\]
timestamp 1644511149
transform 1 0 41860 0 1 52224
box -38 -48 1970 592
use sky130_fd_sc_hd__sdfxtp_1  scan_wrapper_lesson4.scan_flop\[4\]
timestamp 1644511149
transform 1 0 42412 0 -1 53312
box -38 -48 1970 592
use sky130_fd_sc_hd__sdfxtp_1  scan_wrapper_lesson4.scan_flop\[5\]
timestamp 1644511149
transform -1 0 44344 0 -1 55488
box -38 -48 1970 592
use sky130_fd_sc_hd__sdfxtp_1  scan_wrapper_lesson4.scan_flop\[6\]
timestamp 1644511149
transform 1 0 41952 0 1 55488
box -38 -48 1970 592
use sky130_fd_sc_hd__sdfxtp_1  scan_wrapper_lesson4.scan_flop\[7\]
timestamp 1644511149
transform 1 0 42320 0 1 54400
box -38 -48 1970 592
<< labels >>
rlabel metal2 s 7074 0 7186 800 6 active
port 0 nsew signal input
rlabel metal2 s 41206 59200 41318 60000 6 la1_data_in[0]
port 1 nsew signal input
rlabel metal3 s 0 27148 800 27388 6 la1_data_in[10]
port 2 nsew signal input
rlabel metal2 s 57950 59200 58062 60000 6 la1_data_in[11]
port 3 nsew signal input
rlabel metal3 s 59200 49588 60000 49828 6 la1_data_in[12]
port 4 nsew signal input
rlabel metal3 s 59200 36668 60000 36908 6 la1_data_in[13]
port 5 nsew signal input
rlabel metal2 s 50222 0 50334 800 6 la1_data_in[14]
port 6 nsew signal input
rlabel metal2 s 21886 59200 21998 60000 6 la1_data_in[15]
port 7 nsew signal input
rlabel metal2 s 24462 59200 24574 60000 6 la1_data_in[16]
port 8 nsew signal input
rlabel metal3 s 0 22388 800 22628 6 la1_data_in[17]
port 9 nsew signal input
rlabel metal3 s 59200 57068 60000 57308 6 la1_data_in[18]
port 10 nsew signal input
rlabel metal3 s 59200 14228 60000 14468 6 la1_data_in[19]
port 11 nsew signal input
rlabel metal3 s 59200 46868 60000 47108 6 la1_data_in[1]
port 12 nsew signal input
rlabel metal2 s 19310 59200 19422 60000 6 la1_data_in[20]
port 13 nsew signal input
rlabel metal2 s 42494 0 42606 800 6 la1_data_in[21]
port 14 nsew signal input
rlabel metal3 s 0 1988 800 2228 6 la1_data_in[22]
port 15 nsew signal input
rlabel metal3 s 0 57748 800 57988 6 la1_data_in[23]
port 16 nsew signal input
rlabel metal3 s 59200 54348 60000 54588 6 la1_data_in[24]
port 17 nsew signal input
rlabel metal2 s 17378 59200 17490 60000 6 la1_data_in[25]
port 18 nsew signal input
rlabel metal3 s 0 29868 800 30108 6 la1_data_in[26]
port 19 nsew signal input
rlabel metal3 s 0 40068 800 40308 6 la1_data_in[27]
port 20 nsew signal input
rlabel metal3 s 59200 21708 60000 21948 6 la1_data_in[28]
port 21 nsew signal input
rlabel metal2 s 11582 0 11694 800 6 la1_data_in[29]
port 22 nsew signal input
rlabel metal3 s 59200 31908 60000 32148 6 la1_data_in[2]
port 23 nsew signal input
rlabel metal3 s 59200 16268 60000 16508 6 la1_data_in[30]
port 24 nsew signal input
rlabel metal3 s 0 7428 800 7668 6 la1_data_in[31]
port 25 nsew signal input
rlabel metal2 s 23818 0 23930 800 6 la1_data_in[3]
port 26 nsew signal input
rlabel metal3 s 59200 44148 60000 44388 6 la1_data_in[4]
port 27 nsew signal input
rlabel metal2 s 37986 0 38098 800 6 la1_data_in[5]
port 28 nsew signal input
rlabel metal3 s 59200 6748 60000 6988 6 la1_data_in[6]
port 29 nsew signal input
rlabel metal3 s 59200 51628 60000 51868 6 la1_data_in[7]
port 30 nsew signal input
rlabel metal2 s 38630 59200 38742 60000 6 la1_data_in[8]
port 31 nsew signal input
rlabel metal2 s 28970 59200 29082 60000 6 la1_data_in[9]
port 32 nsew signal input
rlabel metal2 s 634 59200 746 60000 6 la1_data_out[0]
port 33 nsew signal bidirectional
rlabel metal2 s 50866 59200 50978 60000 6 la1_data_out[10]
port 34 nsew signal bidirectional
rlabel metal2 s 14158 0 14270 800 6 la1_data_out[11]
port 35 nsew signal bidirectional
rlabel metal2 s 59238 0 59350 800 6 la1_data_out[12]
port 36 nsew signal bidirectional
rlabel metal2 s 54730 0 54842 800 6 la1_data_out[13]
port 37 nsew signal bidirectional
rlabel metal2 s 26394 59200 26506 60000 6 la1_data_out[14]
port 38 nsew signal bidirectional
rlabel metal2 s 34122 59200 34234 60000 6 la1_data_out[15]
port 39 nsew signal bidirectional
rlabel metal2 s 52798 59200 52910 60000 6 la1_data_out[16]
port 40 nsew signal bidirectional
rlabel metal2 s 57306 0 57418 800 6 la1_data_out[17]
port 41 nsew signal bidirectional
rlabel metal3 s 59200 42108 60000 42348 6 la1_data_out[18]
port 42 nsew signal bidirectional
rlabel metal3 s 0 42788 800 43028 6 la1_data_out[19]
port 43 nsew signal bidirectional
rlabel metal2 s 36054 59200 36166 60000 6 la1_data_out[1]
port 44 nsew signal bidirectional
rlabel metal2 s 21242 0 21354 800 6 la1_data_out[20]
port 45 nsew signal bidirectional
rlabel metal3 s 59200 8788 60000 9028 6 la1_data_out[21]
port 46 nsew signal bidirectional
rlabel metal3 s 59200 29188 60000 29428 6 la1_data_out[22]
port 47 nsew signal bidirectional
rlabel metal3 s 0 55028 800 55268 6 la1_data_out[23]
port 48 nsew signal bidirectional
rlabel metal3 s 0 47548 800 47788 6 la1_data_out[24]
port 49 nsew signal bidirectional
rlabel metal3 s 0 44828 800 45068 6 la1_data_out[25]
port 50 nsew signal bidirectional
rlabel metal2 s 45070 0 45182 800 6 la1_data_out[26]
port 51 nsew signal bidirectional
rlabel metal3 s 0 50268 800 50508 6 la1_data_out[27]
port 52 nsew signal bidirectional
rlabel metal2 s 7718 59200 7830 60000 6 la1_data_out[28]
port 53 nsew signal bidirectional
rlabel metal2 s 4498 0 4610 800 6 la1_data_out[29]
port 54 nsew signal bidirectional
rlabel metal2 s 16734 0 16846 800 6 la1_data_out[2]
port 55 nsew signal bidirectional
rlabel metal2 s 52154 0 52266 800 6 la1_data_out[30]
port 56 nsew signal bidirectional
rlabel metal3 s 59200 24428 60000 24668 6 la1_data_out[31]
port 57 nsew signal bidirectional
rlabel metal3 s 59200 11508 60000 11748 6 la1_data_out[3]
port 58 nsew signal bidirectional
rlabel metal3 s 0 9468 800 9708 6 la1_data_out[4]
port 59 nsew signal bidirectional
rlabel metal3 s 0 4708 800 4948 6 la1_data_out[5]
port 60 nsew signal bidirectional
rlabel metal3 s 59200 1308 60000 1548 6 la1_data_out[6]
port 61 nsew signal bidirectional
rlabel metal2 s 9650 59200 9762 60000 6 la1_data_out[7]
port 62 nsew signal bidirectional
rlabel metal3 s 59200 18988 60000 19228 6 la1_data_out[8]
port 63 nsew signal bidirectional
rlabel metal3 s 0 34628 800 34868 6 la1_data_out[9]
port 64 nsew signal bidirectional
rlabel metal2 s 47646 0 47758 800 6 la1_oenb[0]
port 65 nsew signal input
rlabel metal3 s 59200 39388 60000 39628 6 la1_oenb[10]
port 66 nsew signal input
rlabel metal2 s 12226 59200 12338 60000 6 la1_oenb[11]
port 67 nsew signal input
rlabel metal3 s 0 37348 800 37588 6 la1_oenb[12]
port 68 nsew signal input
rlabel metal2 s 28326 0 28438 800 6 la1_oenb[13]
port 69 nsew signal input
rlabel metal2 s -10 0 102 800 6 la1_oenb[14]
port 70 nsew signal input
rlabel metal2 s 35410 0 35522 800 6 la1_oenb[15]
port 71 nsew signal input
rlabel metal3 s 0 12188 800 12428 6 la1_oenb[16]
port 72 nsew signal input
rlabel metal2 s 31546 59200 31658 60000 6 la1_oenb[17]
port 73 nsew signal input
rlabel metal3 s 0 19668 800 19908 6 la1_oenb[18]
port 74 nsew signal input
rlabel metal2 s 2566 59200 2678 60000 6 la1_oenb[19]
port 75 nsew signal input
rlabel metal3 s 0 32588 800 32828 6 la1_oenb[1]
port 76 nsew signal input
rlabel metal2 s 1922 0 2034 800 6 la1_oenb[20]
port 77 nsew signal input
rlabel metal2 s 55374 59200 55486 60000 6 la1_oenb[21]
port 78 nsew signal input
rlabel metal2 s 43138 59200 43250 60000 6 la1_oenb[22]
port 79 nsew signal input
rlabel metal2 s 25750 0 25862 800 6 la1_oenb[23]
port 80 nsew signal input
rlabel metal2 s 59882 59200 59994 60000 6 la1_oenb[24]
port 81 nsew signal input
rlabel metal3 s 59200 4028 60000 4268 6 la1_oenb[25]
port 82 nsew signal input
rlabel metal3 s 0 14908 800 15148 6 la1_oenb[26]
port 83 nsew signal input
rlabel metal3 s 0 25108 800 25348 6 la1_oenb[27]
port 84 nsew signal input
rlabel metal2 s 9006 0 9118 800 6 la1_oenb[28]
port 85 nsew signal input
rlabel metal2 s 18666 0 18778 800 6 la1_oenb[29]
port 86 nsew signal input
rlabel metal2 s 30902 0 31014 800 6 la1_oenb[2]
port 87 nsew signal input
rlabel metal3 s 59200 33948 60000 34188 6 la1_oenb[30]
port 88 nsew signal input
rlabel metal2 s 33478 0 33590 800 6 la1_oenb[31]
port 89 nsew signal input
rlabel metal2 s 48290 59200 48402 60000 6 la1_oenb[3]
port 90 nsew signal input
rlabel metal2 s 45714 59200 45826 60000 6 la1_oenb[4]
port 91 nsew signal input
rlabel metal2 s 5142 59200 5254 60000 6 la1_oenb[5]
port 92 nsew signal input
rlabel metal2 s 14802 59200 14914 60000 6 la1_oenb[6]
port 93 nsew signal input
rlabel metal2 s 40562 0 40674 800 6 la1_oenb[7]
port 94 nsew signal input
rlabel metal3 s 0 16948 800 17188 6 la1_oenb[8]
port 95 nsew signal input
rlabel metal3 s 0 52308 800 52548 6 la1_oenb[9]
port 96 nsew signal input
rlabel metal4 s 4208 2128 4528 57712 6 vccd1
port 97 nsew power input
rlabel metal4 s 34928 2128 35248 57712 6 vccd1
port 97 nsew power input
rlabel metal4 s 19568 2128 19888 57712 6 vssd1
port 98 nsew ground input
rlabel metal4 s 50288 2128 50608 57712 6 vssd1
port 98 nsew ground input
rlabel metal3 s 59200 26468 60000 26708 6 wb_clk_i
port 99 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 60000 60000
<< end >>
